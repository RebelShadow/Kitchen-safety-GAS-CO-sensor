PK   ?T$�2@'  �~    cirkitFile.json�ߎ�F��_Ũ��US��$ug{l����c�s.,� ���X�K��z<�t^�<��`uK]d����b�F�����Kf?l��ߺ�j��w�ߺ����n����z��V?���ټ������}������sv���.k�]�6�Ԧjmٗ�n2W6.��2��ES���e�U�2��?�����-���R��b�S91�Ԃ���Aj�TA� �`�(f`��ow����uw�*����e�Ql(�~Ssk2cͶ>�o+�62�\�/�`�B� �`�R� ���<ɊM$
@����.{��<l3jc���۬p�ed�os��u�����9Zl"Qȳ��D���i��D!��b�B���&�<�M$
y��H�+6��t�+6�(�r�~�,i����3 ��y����`Ⓛ��ߺ}��o�-7P�߽����dw���癕�p��D!��b�B���&�<��M$
y�H�.6�$�<��M$
y�Yl"Q���D� �R8�#��]'ϻb�B�w�&�<�M$
y�L\S�4��9[l"Q�s�؄��<g�M$
y��H�-6�(�9[l"Q Ɩ�y����D���]��D!ϻb�B�;�&�<w�M�*�D�D}���y$=#n:��H���&��]J�(��@l"Q ^6�A�8�H�ǁ�D�(�	���@��%��3*�)P����.��D��ˆ�xt�	ȟ$k��T��Ǫ�M鮾�~#9���$��PLE�KF�K�#,��,�w�;(a�L尾sX�A�K�&�w�;(a�R
뻀����t����]��JGX:S�X��X�A�Kg���;(a�LUb}Wb}�#,϶w����Gg���E3t�T��u	Z���	X�X�X�`���s���,��xV9�`���#0χ�,T�|���`���
���|��?�`����WO��-X>�������G`>^��K,��x��`���#0����r�v�?,X�����?�|�W٣5�W�,_,X�`���K����,��x�`���#0/��,_�|�ㅃ`������|���?�|����k��������|���?�|����Ȃ��/X>���^��������OX8�������D���X>��bn�����G`>^��X`��ǋ����,��x�>�`���#0��σ����|\2�?�������=���X>�q�
�����G`>.��z�	z�	Xx���`���#05��?�|��r,`������|\H�?������K����X>�I��=�:���_U��q?X�����/S>��$�� V?�~�|��N`������|\O
�?������+a���^e�^fV?�~X�`��������,��̤���>Qw���>��)��Ӹ���`�4�]�R���`����G`>���X<a��ǥ����,]�[Yo\
rm9=Y�qŕ�ǕpWW%��}���J�qە��wi�|[w>p;�y[��)�͊�L��3��#+�<��EG&ɑ�c/��^J�Nr��')׶޶�o9�m/�q'�O\�^x�M�Y��),��E�X^�~\�x�@ʣo�]��@��w��x�|�Xrt�}4���������B�\�>�3h�����[o�u���_z��q�]抮�|۬�y��>�L߷1Z�b�sA����e�m��7�\V���ΣuT�ν��]�������d}���'#Yi�2��oLM�mQ�x����5���[��c�)o��r�b[�m�l���/}Q���/,u'{����	Pd����ބؖ}�gul��G�fM����2���Ml��aQ��˰����kQ��.�B�!(�>��[�:G�{^�6/��4YW4u�o�t��L����mx�_�|�޿�î�������$��D��3���Hn����`�@��'"�!÷�d��H
�d���
�d�� �h0��ƭ�(G��������a��"qY��-�m�L�č�d��/,w,y�,�a����K�(KfH1�r8��8ʒF)AL�<nayeiM�ʐ���B&\����q��O�� f��q�%3��`y���8ʒ�AL�<naye�C� &Xw�<��d��y,�;XGY�2I0������2��8���1���q�%.;c:Z���5	�`ye�ˣ��`y���8���1���q�%.7c���ay���8���1���q�%^c��q��(K���'&g
�<�F��*�>Z0��8��0-�ǟ:c�N�����Q�x�'�	��,��,�BD,����`y<������GY�%2&�B&X��<>gi���;��a���d��{S<C��ݵ��x����a���J*���Ѓ[�U��TXM5�[�
��+��&ݥ��qU�4XI�5��T�:�v��+���>��_�UP0�`%VS�������J*���K�[�U��TXM5.��
��+����%QHa���Th���P�KIt)�.%٥��HGx���R�%Z�k��[��BK:�<g^Ƿ:
L��thyouT�
-�����(1Zҡ�:��Qc*��C�kJt|���ThI������VG��В-���y����ThI���*��VG��В-�����1�Wb:����2���Th�<�|����2���ThI������VG��В-�I��.S�%Z^[��[]�BK:��FTǷ:�L��thy���out�
-���]��I:�L��thy�out�
-���j���2Zҡ��:�U���4]Q�}���eNG��В-����.S�%Z�1��[]�BK:�\+AǷ:�L��th�惎out�
-��r�
���2Zҡ�*��:�L��th����out�
-��rM���2Zҡ��.:���e*��C�5jt|���Li)��.�:����2Zҡ�A:���e*��C˵�t|���ThI��k8��VG��В-ע��.S�%Z����۠����"Jz��rm0���2Z:O+�ttY��e*��C˵�t|���ThI��k���VG��В-����R��2:�,�負��ThI��k��VG��В-�d��.;C���負�˂�.S�����m��eQG��В-����.S�%Z�Y��[]�BK�hW~�z���J+3�iWZ��&���L�V����J+3��W�|�B�{���uI0�~#�r� =�g���P�yZ�}mԁ��s}]k�s�V]k�s0]k&?�Zkf��Z33���f=L�}�s�L�R9���Z3�(���Z3�(�3_�Zk�� �ȭ5���O�5� �q�]抮�|۬�y��>�L߷1Z��W���E����]���`+���c�ɵ��ܹ=�EV����d}���'[Yi�2��oLM�mQ,aY`�"K�P�Rm���1�YI9e����m�}���,��\d){��<l3jc�nY�+����y��>���e�����̗�?YiBl˾�:6]�o��O�gc���&6��_Y��EV.>Y�أIN�֝�L�m��MimV䔼��hԙ'����Y�K����e_�&늦NQץ��k��2�魯۰�>Zb��5�}0Sv���>t��>�]�������s��_� :�B2d�؆���>���AC�@�̠�!D CfP�"�!3(}ȐF D Cf�����h&E�6.m��6�7ʒ9�`�`��`�e���0L��M���d�]&X'XGY2�!8,�[XGY2��A�������q�%s�0���q�%s��0���q�%s7�0���q�%s���qXw�<��ĵ�`L���P
,�;XGY�=0&Xw�<���5b`L�<�`ye�k���`y���8����1���q�%�� c���ay���8����1���q�%^�c��q��(K������,��,�ZS,�XGYⵍ0&��M��MX�<���k�`L�<`ye��<��`y<��8����1��x���9K���L�c���� ��
+���j�m�WVRa5�d�*Я���j�Im�U�_5XI�5�.�N�b@<��J*�����II�4XI�5�QT�:)��+���jRm�WVRa5դ�*Я���j�I�U�_5XI����ťBK:�<�YǷJ�KIv��.�^���ThI�����VG}�В-ϙ��S�%Z����[�BK:���AǷ:JL��thy-��ouԘ
-�����(2Zҡ�1:��Qe*��C�k|t^,��2Zҡ�J:���e*��C�k�t|��FL镘�.�:����2Zҡ�5p:���e*��C�k�t|���ThI���$��VG��В-����.S�%Z^#��[]�BK:���UǷ:�L��thyͮ��$]�BK:���XǷ:�L��thy��out�
-���Zp�*�VT����˜�.s:�L��thym��out�
-��r����2Zҡ�Z	:���e*��C�5t|���ThI��kW��VG��В-��P���e*��C˵Dt|���ThI��k���VG��В-�v��.S�%Z�Q��[��dJK�tt���e^G��В-���.S�%Z�}��[]�BK:�\�IǷ:�L��th���out�
-��rM-�]�BK:�\LǷ:�L��th�ƙ�out�
-��r�6���2Zҡ�s:���e*��C˵�t|�T�C�̇�.:�,��2Zҡ�Z�:���e*��C�5u|���ThI��kK��VG��В-��T�m��e*��C˵>u|���ThI��k���VG����2�矢��/��bC��꘬Z�k�m�p~;��VfjӮ�2SMv���:�+��T�^ie�V�J+3խWZ��G���L�Vfj>��:P�b�wk�`�w�Ӫk�`"x��k�`bx�3�k�`�x�c�k̀r0&��R��&����&�羸��&��k�����⹯>7S�m^t�+�2�El�"�MV��3}��hݒ^�+Y�2�6wy�Ƃ�t.�C�YL'�:*s���YY�����M�3�le��ˬ���15m�E��e���,]CaK��
���S�f%�Ŷ�۶����/�,�r���)��ͨ�ɻe����.#S�}��<���,��\diBl˾�:6]�o��O�gc���&6�2�"+���EV.>��u�g�y��ySZ�9��5�Qg.�e������˾(M�M���K��63e,l�[_�a�}���s��o��~���w�}u��}��f����޿��][��U�}��7��I lDt4"���z�ԛC��>A��+;�1V)N�?�DiF�3�HkJ�N�KA�@5��."�ỳ�����а����2�%<�u�XWU���d��X�4I����n����$c��#K���֧��/��U��B�"���e�߾}�g�_wK���=���)A1Ϸ#B�?�}�P�7
��vJ1��M1�.*�
�S}��翧�~�<�Bڏ�o�k�\�"��: �F,>�=
�>��#�3�q���_!�� B����l_ʿ�U�~�[��nI�j~��<��s����ݮ�?ԇn���ϻ�?�:쪇�v����ǯ�����/������Bl��&�bfx�)��0�dE!�؄&;
)�&�0YRH�&�ɟ���*�C�M�aBl�s?�b�8wT����Mi�A�H�r�8V�ȰH�r�8W�ȲH�r�8#X�H�ȭr�8'Y�H��^�6�qV�(5Z!���ҫ������$�d[�s�7.� d[ȶr�8s]�ȶ�m�6�q�m ��m���}) �:@z���O9 8��ՔB,@z���/ 8 ��ҫ�W�p��p)�X�l+����l��Vn�i8 �����hp Fcñ����Un���8 ��ҫ�_p ��S��a��䑕˰ ���Ё�B,@��l+�1�{��G4�LG�R,@����~ @���+��U� ���i�
 �r��X��]]��a���=^������6֗���I��;֙ٛ�ݘ\J᜜	�Ⱥhr��&�҄ޝTHz�G`>SM����A���#0��&��q� ����/���&U����#0_ꛀ�7�$-<_,��R/�I�h��b��g�Iah�=���|�3դ�3��X>�jR�g�?,���ɔyL�O���U�	2Q��&���*A�B�B0!�	yz.ڇhq&$4!O-F�-P���&�i�h�E
��Є<��C�P�����}�+`BB�Tz�тLHhB^��!Z��		M�K���h�&$4!/�@��S���&�"h�_��ߠ�u�E�q	�)�uʔp4!|+jѲŢe��Є���C�l���F�}��-`BB�.�ѲLHhB^���!Z��		M����>D�0!�	y- z�Z��		M���>D�0!�	y&ڇh�&$4!�E�>�>��zšu�C�0!�	y�.ڇh�&$4!/2F��S���&��h�u
��Є���C�N��W��}��)`BB�*z�=Z��		M� �>D�0!�	�zڇh�&$4!W^@��S���&�h�ש���u�G���)`BBr���:LHhB�4��!Z��		M�UR�>D�0!�	��ڇh�&$4��|�j�����z�w����ks��e�p����+]���	h&$4!W4B��b���&��Kh�U��Є\:
�C��{��{��	h�*LHhB.م�!Zŀ		Mh&�c���pB�Ru4�}�KѢf�qj�KѢfJ�R����h��LHhB.Q��!ZԀ		M����>D�0!]"\���I�ŕ�'5�~�S�~R ve{?M��/�N꯮���dՍ�3�������TB��;S�4HBQ��`�~�n�i8O��ր4���h[k���($ߤ�~$m��IYܵ9N��I����B 7}0Z��of�5 [{�3*k�I��Ğ4���{Zk���Z�m^t�+�2�El�"�MV��3}��h��}��_8~]��.��Xp��eu�1��TZGe�܋}�E�_<��nkL�7��|����/�����Դ����_����w�-�&+\3Oy���S��o�f���~���ڿp��b�*�Js�����\b[�m�ձ�2}�5}
1�P�.6��/ygQ�����9}Q���kۺ��l�y��sSZ�9��5�Qg�]����"sg��L_��y��ɺ��S�u)
��f���mz��6�x�,i�:��l>��m�îJ����Y�7���c��3��f��Iq�q$�kW~fp���Ò��Q?�r���C��O܀���v��-,����r�-,����r�-RZ~{�i�Κ:�O�w�����>�k�ƾ���e�'��fj���hR0��quWvY��4�_Eޕ�璤��%���,:jp9�4X��N,�$'��k�8H���'� n�5H��pٻ��[�Ҩ�1�z5-��M�HG�Y��)�=���K#Ё�)���B����0J�bq(H]&�)� E)����tbʔ0�
��1��4%,D��73EJqJTJ�$af�>��Ȋ^1M�M	���Jr��3Dn����-7��x	��5g�di��9�����f����)P��\���^W�Y<t?T��{�}�Q�bU����+>�h=n��&���N7��Mn��?n��M�qS�n����tS��)�n*7�M��r��>������iz��t�4=kz:k��6=�6Mϛ��M/=�$�']��ݻ�Y�����������qQ�DW��/��H���r�UF��:=��]���Y���κ�C}`��a�����n��5���;��o���������Ȼ�W����l�V�{����D����t����_v�����dw���wi�}�����m����}�n�]�y}Hg�.Ư��C_o�n���ݞ��ۇۻ�$������v���S���UR��7��B�&�1��X�6���!�,�f���6YѸ��<��s������͢1���n�.W}��<�O���������7�4oo�gg6�\3�"3-b>�"̵�s-hfC(gL�b�E�k�Z�����ō3a�U_��?���G��6x��`�Z�L�Xδ��\�8�brA�6رO�6L����z�0�RO&W�i��J=m�\)��v�-�����᡽������ze^ٔ��$���ܥ��,�@�fO������+�HTPH'���߶��L�Ӿ����N}H�,�6ε&4�����_4�8����?�r����M]�W��>�\JP鹘N׽*B�bJV�9O2\S6!�q�..u��-eu�R������ЌOw�`��t�'�l7����a�=K��'��ϒg;}z�<{����;z��b��Z޶�Q�����dn�Կ�����GAY�(��{���4	���v����^�p¿��޳�!�Wv��yE�����[�����W~ޟy N����k���s��7�]{�"�x�g�'��&��E�?�J��tcG��On��n�6Ĭ�k���)s�!����1�-���>y�/��)n~c��K���G�d��_�����ü���0l�Y`/z��(��eq}f�qX_�k$������!sy�_��f���t:pB>�*˿�?��:���?�*>�M�@-e)�z���X�Yߛ��v� �G����8|o��y�&/}��i�xn�F"�
� Z�yQ M���ɿ��ܕ_@�|����������n���Cl��@�	����Mf����A_�R�[\鲦܆�hL�m�o�t�k]���;	�E����$/�#:����:���Ȝ���~����?�)��~����b����_}�ql6E���&|�7n*>޻���,��Qt}jص�u���<s���Ge�͢�'��R`��ˍs�Y�8�Lv���nd��;��Ğ~.sË����%�����"���~7���<yW���G�6�m\
(�c]�Y���;�Cݥ�4��E���(:�&��i�v�aHi��_7,v�����SR~&I����If�D��b��d�ݒpv6?Mvgaҗ�����m��t�vɡ��m�+�)�۠����������n��/l"��*F����K7�Ŧ��+�������m�qz �7[o��o>���a����m���Nt��oҝ�n��y�f�/�϶�lnޤ�Y�?����6]=;q0�ݵgLI'+���o?"Q����h��n�?ԇ_�޼y��7���?O�{������ا@�����{ܜ�-�pv��W�b7��}�����)�N�'�Ѐʵ���=��:��6|���+���>��&�nùݞ7_�-���n�lA��f04�F��/E�'�������W��g�s�+�Ο<>+W��Z���i�I�� (W�A �
p~m �|I ī2������ X;�]�zG�t��b]{y�E�w�W<��k��a�D��ݦ���Wv�:�8\����Ɓ��&�\�$��{��*������f ��mi��<�^�x�%*��x1b�׆�_����l �� 0
 ���-���Z�����5A�WT�=6׺��׵���������XY�~/g����d��.��ɳp���\~�.�O`�Ȫ�ɇ�a���Ny�$:G;��n�i�g�nK�E�7�+���BH���9��9��#�KR�h����2�q_�{3(�-��^l�>�lAW]�������W����t7{�|&��p�n3ͼe���h��i���_g,[l��и���
4TH��R�iD���S�Wx��m���|�����>�Uh��~U�zr�?�"�����^�ۙ��gzq��5m�ZG�����gh� �
ֵQeG���Ib�M����ua�|�#����.pDw_�U�t&��m�_��iX<��_�p��~I\�}�Wv_V��XV������+X�����G/���eoE����PK   /�>T�a��V _ /   images/b9b5db0f-1139-4dc1-aec6-3976f40bff5b.png�S{%\��;3c�۶�b۶��m�b۶m'��̠b�o�}������O{Fo���SQ
   �H��  @  ��?b`B  d�EԼ�>-�7�J���Åo:���bfb1��hEAh9vU�p]��ؖ-L9ǈ>��4s�c%�3˜m|68�A��U]p���*�Sbk��O�A�kWCq 䊙:�b�6·C����,�yn˶�Z��E�8V'�h1������������52�?p�"U�L?�_��	*��l)Γ�Z���Yw{L����׎;�${	O
j���
�?;�xW��R}^f��^��PB
�ز��~�&�o�s��k7͵��v%�=�����������Ѣ$��鷢$M����O/�q���Jx�+W�s�ܘ�bj��Y���<t��,��'�ƽD3��4�%O*b@��P�t�]��;��p����HJ��N!hT���A	�?��	���j�ؼy#Q��u�p)n�MY`��L4P(���1^oMBSB>E���*~c�D����!��GR�qHP��$�b
�j��:���yի�m[wfM��|�}{{{����9�.�g�R��Q��gb�[��8����������#�6~z�33K�D��~��Q���@�7h�?C�_Ǩ�[q����Of:�$��(���~��x)��?⤂Xr-���I�O-��1T����>4���?F9 �t��Zw��ڎ^S&�JG)�;/������*2%G�gg��q��]������͋n�Z���;s���vv3|3�uu:�� �ǒ�Ic�mw�6ݵO�M�a���}̳aLǹJ��b���K��:"�A��lɛ\��������`�O�����ےb=�3�V�e�5} #n@���Nq����4���P��G9 ~�6��	 �J`ͤY���1T���a�+Uq���e\O���a���P�i8�۱���ɘ��M���+/F95o��}��U���l~ʥӬ�Y�-_fL�ꪬ�ѤƸ�ŋ���"�˘���Ȉ.�z�����S�ZrXm�0.e}�F���gu���7��JT��h��G����n����!���0b�԰r\��5r��<�c���(�s��j0��!�p�����{Iql�sRlpOf��R�n&� �Y��>(K����l���γ]���*�׃�(l{k�E�Y��f)n0�?����v��#2���;.�8��� ՟9���ݎ�a@j�^�`r ������	�P�}���:T���}R-�T8S�8���ۅ{A� �|=�qE.��ta
�u��ۍ5��'!�J~�:F�"�O$�C���+}�F����R�<>Y�������T|$|��c��0�{���r|������fb7rgg�=_�����Y JU�ڍ���VWlm��&2	%eTM�>�t��D/0�
���,y�~��dHS���T�fZ�aBގ��	���*�ߍ�yX{<�A[D���a^t����n�%X6�Ӡ��6b�I��w�,A���-<�s�+�\B�F�g�y���u��3^v	�D{�:��B������,G"���K�%��cfkq�y%�7�����=���^��'������(��"UR��o�tKwu����-�Z�����]ǜ��`i�5pdK�2�H��(��ª?�������#�L��K|�ڍb= 2��0�r���48���M�Pw\��JİXc{b7������U�=��}�u]1�� iA
�FSTtWS�:Nj&�����^���l�zWu�p�������W�IӒ�mK��˼���F;�/=y�&��Dٱ��ef]b�j��~���m�����k�l�ߢJ���PǨN.f�&-̟m���:s�z�Й��6F�*~���Z��\����^뺂h�P���W���)�"�H�ʗ�{S�� N�3�4kT�p%az R��괋�8�8V��.'y������K�D� ���q�j.����8��߸�G9uz��'"�B�V�*A�-|��l:u0���l���k��3���j��ԯ�u�|s �,�$-E"8�������GLKe3�Qi�c��d�a�U�'I9h�X�m;��������O:�9��ݙ@c�v�5�e�e�o5NS������Պ\����������-pb�A�!K� ��<rS�U��W��It5g��ZܨqT��sۤ�O�5��"��rŭ�U[�����NSo_֧��k9�(�I 7ZOĤ�����7S�$����>��t��d��,x"yn�#�̓����py�.�4PP}���^���m���j�����#ʻ
�BY�>�SkK������S�4�7�Ws-b0*0v��pptfu�~�k��"��\E>�����)���c�ԇ�ZV{;�!ٷQ��������m�7���	��V&�Y������E�}kdI%	CR��	}�H�H߅��Þ':d���+��K�I_�=n��q�����F~NY0! vin[�g��cC� Q��\-)���9@�z@��Y��XB��;MvVE�Ǳ�`j��{�1bv�N�y��	��z�o_{4 u�h�e�����3�_�T�#�E���ؤq��_�3�&8���0�y��(��y�G����z��)r�W�YH�Ȱ��A-�Z��wL���3�p�u35��Sq܊8�6�,��g�qJd�u)?ɜ�)l#Uy�.����""�N��xd*�ϊ͑��ޡ�=�4O$�78��� FIR�W����[�>v��� vwt&��6f@�ѺI3�.����kB�h3��yݘ��:,k���
Ɔɘ����xP5P��
XYP��/`m�&P���;��0���i}jI;g��.�L�ฐnIJ�SD�CU����J���hޒ�"���/�4�I>kp׵*^3:Q�	5�_D/^u_�����ަ&�^�r;��6� ����Z�/e9�.CO�w��B�a'-��۪3/Y�8n�}�^����W'��,ݪ�Ŧ�p�����Ǐ@G'��a��co�ݰeLz�)?�RԐ79~�d���,I�v�U|�zt��s�ܵZKc	>�8��ۿ�;��ֿ)5[<i������Q��T�c�Y9[o�~�Oӿ�k�t:�~\�l�pq��I�;p���o6a�@j
� �|���'ڥ��B��E<�h�W��MM|��R�֋fqI�ՊI���Y�?�Ҧ��UG�E>�u�q ����F&���m�V����(��̿=����l����(�R�kC��h��Zh����3)�j=���y(�2�Y�DξK���AD�.��%^�q+�'Z�};_�[�f��1̝=vU���N�V��ښ�,�f;�9�|r��j���݌0�u�xn����`Z��Cˑ�!��(�!�D�k�5&B��W�>~c��Y��-���L��0`�K��5֘F���6�����ƚ1�<ПP\A�&�w���Ex��������eL��.��r�3�<�~s)H!0e?̖��P���
�n|�nP�D��y�آ�0�立 W�`���g	3O{����l)bd�����%�d���<9�������Ԇ�
�Y�$�S�������Lb� O"̣����!���PP�Ey6m��~k��p��q�������y���Y�*Q�М�:��G@��؆�j+3{/�
�)~k/꡸�thf��=F��`��5�)��g� b���7�e�y��M;�}�F�jM�7�,��DOSi�*��3x���/�?��$N�*;9Nކ�k@4���=��lE�KzZn�u0��c����0�f�k`�X(��H$
f�9Y������)�K�F%��oP�-� n�Y�_m5�AK��췊��|%�#v~ �����IE��;����Pp��H^��\/d,������$�����O""O)�َ�}�a-�,T&0���ԟi+��W@Ukᙇ�Ak\�Tp#��8|1q\�Up�p������I'z��� c�0Ҡ��%+5SM�n�f��T��b5�<v�u��'H^Bx�ʹ!�-��1p��?��l#[�XT�z����I�$�3��3�U<LR����E���Q����n��{�eჽ�Ԥ鄑ϑλ��S�1<�Q��x�ì[�t6�R�;�)�������Ɯ:k�^q�E��i��E���i�8���{:v����~�gG��D��kUT�*W���q�qĘyP�k��z�0��� �ӂ�q�*E�����#FI�BdfQ�ڡ�I0���/���aZ�l�� Z�4[#)��DM	��P=�b��.I�J�l]�om��t�YT /�l�2K��� 1�����P�W$��� ��/���Ʊ��6���6��)�o�l�[�P��O��RI���;^��x��FnW�l�Y��Y?7�t'�]5�+7b=K*�FηF��_Pnd�o��'H{��[���ϏsyWƴ&g�I���3���Ud�E�:�dd��������� ��H�v�"�? Σt�;*[cu����/��Ύ�]f�F��ȯ�}���3V�w�cDQ�-�tWY	S�g��O]��n�H��FS<e~�+Tڎ��De\�걡M��*; �a`&\jzR�y�o�Z�*�9y���2G�[f�[��Ĩ�S",����U�*��
�Ǚ��+��3�����|��7lFw��k!��!��� ����Dl�@T�x�.�]QL)P޽����l��9D���^�N��` ��#i�G$3���g�����_��F�C>��p�r�XnE�<��]<ɵWf"ۚ�ڳ����
�*0�BĴy�g_q���t"�D��iу{��kӊ�#�����A���H��m�*3f�G���M�>�z�
W]��s���=x�|����M*d�T�����2Ae[�&��"
]��`NU�K^ȵ���:��M6���4N��5P;�\��/�4x% %8}̝@���d�Xw_�	H��/$����k��Gi36�(G<G�@�/e������ԡ���Ppc�;DAF�i�)hr��#���o�����En�rt)�H�)R<O"|	�}>� 2 I�`�.�&�en�k��f�Q[h(0K
-�لtv�ЪҪ�����_���
%���I�t�Qg{u�%B'>F�n5�������,ꦹvuLdX7�\�{�F����)��яs�5{�d�Z�s{�0�æ��l�O[W�5]�Iqľ�"3�X��ˬ\��6��j���^�5O�U_���0�:0,�+R�*םt!>���?���\�4�qi�[��u�羫�w���%ۍ�Ae;�pڶ��@ep��-�������Ka�����dI��+^
̣���	*T�֧\�����VRG)��>��σ|�ó�����x�^+]T
�!��>��		��.e��/~`̐�e����|[��?i�$EMQ��B���k�jCO��e�Qڽ��{ʏ�;}�]���������Sμ�x���1Aݳ*�����{.@J�b�����|�L�u\Q�:V�,�E`����(N�#�Oö�(�]�������F��O�n%�Xu�u�Z[GxJ����I�b��q����������U���z/G��߻�?�K��~���V%�u�ԫ�*�kQs�Ė�6O��$��F�p�d>�ok��PU�!v���8!i�qx�����vX`LbB� ��Td�฾�J��H��Ȝ�n��� 2W��n��[7WkH���
}P]��x��8�]|`��	���NL�����9���M���6U8J=^�� �G�/���M��V�J���ph[�S2o/�Ӏ���.*��npU�\hx��B!,>7ږl#Hs�b�h���<����M& J�>���/vر#[\��}O��rWe"�[3Z�7 �ƍ���#1��8��p�,Gѱʡ\��y���> ;��vr*�h�&����[d�����ڽ׾�׈.�Aa�C�)�B��g��m*֑�V��j�M{TgwYPQ�Rv�*˵�s�)���m*}~���}�7U�gѓ47*�xY�m�K��Ŏ<�ब�8������4�$?�~�aid�v�ƍs�K��Sq�;�p��s�Y4]������\��&EF�uK|�q�Ig�c4wj��P�}��FdZ��h��U��8	m�x0�|n�!�G�v�n�u8��\��c�Z��=!.�h�mI�)�qD7��"��E�P#�VG(q�C�#W�~b�s�����T3� ��� H�{�p��]�=������6�a�[��a�������ab��W�W]��Χ�(;­�aRا.R�~����y�SlNb	=:_�]��e�e.v��Z����8~}�cJ�)�=��ć�b�7?�GM|���7���;&\��T�%n��G�X"N�©O�S1�	m�����[�8��ն�I:Fw��+��o�'����q�´z�/`S|,�|7���!��gB�=y��p1�Ǻ�E�g�O�fɟ��.m�`A�f�V���m���L6�6"�mň�n�ƕķ��>���6.(�f��n+� ������YN�ы��B����sb��X��Y�*=S��;��v�ر1�I�r��못V@#�hO����PҮP�#dJ����g\��?����4��ԏƿ��0W�X=Z�#,�U̟#}"϶Ly.�>_1�|�Set�u�?R�H�_�
��'3{�/�}����4�;2�k��E�vj��F,�aG��Z�A��l�%��c�
.������F�NR�!�)���"�n��Tv���_$���ep�Q�&�����[e��ِ��)�0��{�}��h�<�ߧt��L� �f0��^ٸ�vd�%�-Q���R:��2�wڋ@;7?�l=��&�je-\ğ4�G�,�+w�����r�Ȝ�:��񀄼yX^2d�1V�p��f �l�9��o��������ftɹ�AM#�@�S&�����C,�yr�˨7��	s�������������C9:Sr��3bc%o ���S#j�����Nl>6���̖��}�l仮������AĹ��d�M��ډC�ۄ!d1vƽ�U�Z���߰i?|HW�L(�1:�aG"�C�V������w�Σ���EL��y�!�_sK7UtppOP\Ӷ�s���lܯ��lPf���y++�Lb���V�Gǵ萢�0�L@�j��8�)C���#�t�5�����F@9"AZ&ѵ�H�W��7���rf^Ji}�5��k��l�Q:y�>Q��k�;�K�i�ɟ�u��}䐈�\a��`�ef�B��3tիJ���y���kZOQ�C����	����B��(�_YD�~d��5.[!�U ��;:��C� @�95-Wa/4O���HAS�)C�՚�u��b�8=�d]e�C#Ǿ(�~w�R����=���x�y8�zgg�+�P�#֛kw�����DIbWrwϳ$^m4����I�y�Fw�o��/�6,T�ld�0�i�vK��x �="XUPݱo!2G�h\<�Ʌ�(Y	r�f�$ѳ�3�L���6�2�>o��ϝѮ��Z��	3�}�bs�.|K���M�.C�+@���[�ۯ��8���w{��Y�R`v��et����I�f��B4Q�T->�I_�
���e�Rx�����-aY4&E��і�C8 ����ğٯ�!�L�," <�v�NװSy�g�/H�t�����_o�� �+U�ht>_�o.}��t���-[���&<2˴�t|+�ms��͂�vB ;��Ph�=B��d����c2J`�t���T[׉pV�R_g��\Q �{�]�B�N'�u[���:p�QJ;{�0������鱊�.�Ą�$�,�2��0���	/E������iV��}��ќמּđf�������0݈����;P1�|["�g�l,��1^:d�T�6�x�A��L������ׁ�pY�/L�>�&Rd �/�	���UKF�棧��`�Ho$�S���R�r7ǞH1ʫ�������5a�@6��Q}��
�B��W����M
: �k�P���1���w�m5��F�Q�4l����e]�݈����T%�M�������(�� ��r�<���
�(�o�m���K�K8����s��p4�I��}�Ԝ���o�9�Q&�A���L��=t��3��~o��?��i���vۻI_k��S=�K����*��Ma�׭e�|C���Q���9���J���U�ۼG����$�Pg"�Đ�eX��r���t_�����=�)n�G���L� ����%Ǆ�O%��`uQw����c����SD�w�؁8:����L����Qȵ�b� &�r)��>ҿ���Bo}p
�(�\Q��֑*N-45����rXT�!�<58������\G\*��4�8��d��nؿ�u:�ѳ5^fxnu�!87}�$ rr)kᠭ�%d �u��
E��+�_��Š���^�[��9�$���`�,�2#���19��r��L3�ζjf�2���<>F�/���{G��&f-F��g^�Y!�W�xN���Ȏm�T�c!labd�fr)pb�b2�+B���o��
5���u|����鑑z=F�Pw��@t�B�o��4�����v��V.\AG`�
��vSJ��g��(���#���u��A!�d%�薗V�|���8�X��9k�r��d�-�����h�V��r���q���ڿU��{���ѩN��<�zt1�c��WK ��6��n��^o���\�@�)
��=�%��Z]�;�R��x������-�}f���l?`�� TΡz�A�"&љC�U �������L�n����6�R̽;�rEqҗ8��vb�+Q��~�?��ZDpr���Xg��1�(}p�����������nJ+֮�":��=�
c��|�9�ry��5�ZV��Q��j� �9 �k,�v�`��������߱B���`���z�\%@0;Ru-���;R��ř؇.�c�TP����.y3�R꾿�Wlz�Yk&Vp)�i �%�u�eC`#*,A �w�x��m6��]r�m*�hp�72��iմ���� )�I�C�*��e�فFRҿi7?�����zZ9)�$���N�4����Ԫ���<���t4��+"v��t5�ќ)�]u���K�N�F\v܄����*nV��V�R���T;#��c�f���v��F=e�f������Q��"陝-	'd$q�"BH�*�1sΜ	�nH~�4?�qf`��4�H��e-M�U�B8k���������HҞW��2%��Ak/A<B�*^ �a�	�]�=�v�NO2���J:�btM�����_��r����IkU\3�N�T�M!���I%Үǀt���Z}�ea��}��^P����fA���Ē�����5�ܢ&*�B�]��\g�\�{��N[4U��2�`�����Z���7[g�70)NrR�S15�M����#R,��,�ڵg��$��nˊ��=MdAT����`�����.�;@h��[<��ܐ�c^)��/Sۂ��D��9Q>CC���&u(���g^�����l���������&4��w�~	�b�<�[~{�N�ݺxi�$��U^1Hxf�m ��VX���Ay��� mC9�U�<�"�kǅ�Rz�0SԺ�����lJ��WN	~��u���i"��CK���Vw"�#��o���w�;��&س�>�ױ���j�yG4�&hW��P�K����7Ab���Q>�]�����E�VãD���
�_#�c�o	,�h�U6I�0*���-8܇B,YW�h�zpQNa3��a|[�z6���CJ~��'�
X;����a�ϳh��7��{n�����.�|�ş�m�����U��Rj?�����jl���(�����WQ0�b�� b:��Z���;ԫ����G�z�mY��z5v�=����<zW�F6qЧ,�y�;��}�?;�
,m�0�����j˴$�Y�� �U�%��:�(0j�D��*3],S[3�c1���O�P��x5m�A�*�̑0'1&%�k�3x��MpV���}w���=�B"p����� ��]�"b0�	�c��[5� �_���k�vs��Lɑ��ء؅��K,Y�j"b`6͍��\�g�s��&T�m7?��JN��wN"x�m��>�1w�;`��� _~�W�be�*5.7M�%���)�~v%�y	��$�w�xwev���+A��;k�L����T��Jk�zjs&���n��c�������� 0`��%q��)�1�1���$pa���ր�MSW�i�B�Fp�V�{Fh7R��3N�w�h�cvr̳��U�S�>b�NV?$�+"�'L5s,R��]*�N�3���G�ȶ��:�7��b_�~�{|��5��\ׇ|�`rxJ ��l|P�-C���|ɡ7�_���
��2I�m�Ќ��
\�v��~��70e�x�rJ
����!��[�y��ۃ;Z � �$h�����/h:�̫�|"?'&�O㺭ZO���ؤ��2�N~�S٪�[i�Tۥ�U1k��7�z#�P�^�oKV�^�3T��x�n�C_��ʚ볎�w����cP�<����T���]�j�;|��%Vu2�cZ�"{V�fRְ~x���q�.�V���D/E�T&GĔ�w�a��-�q �y���~�%� a��r��j�����~˟Y��V��c�4T�����1|�P���8�,9���2媫��H�	r���=t�Y��^\�8ΰ�C}_��^�h}0N�h:z8�/wx�7��+L�'ȸ�`�g�8�{�e����e��%���5s?5]�U�rǂ�X���~�;��q���z�D���G������7'%.��-���xɼ�y�;�A�YA�n��BҖ"b_��ٮ=}a��ڞ}?;#"j��ZC�i_e��$��
�{��EP  �f���[ZC�o�؃�������m��.��Fv�Z�E/����y2�+���S�.G��<��w]�bƯ�Q��8�I9Vcj��W�(+Ǡ���g�����ȇ&�c�}8�ǆfih3>����Jy�C^/ƕ�^�_�vPGg-�@ş��)���'��2��P�!�ە�&��AN?JN��Ү�L��3st��x���#?�2`C����YW����6!���"LY�X$��b���
+3a2�0��p�خL��a�Q��N��UO.�QR�G��F髚��훞�s�ݎ�Yuϵ�7|�z~����76��R\+r�*x�f�UAx������lcu%����Q��:E�E�dS�}R듾�P��g�Ξm���#bI�� ˔���M��7R���k7��l���H��no�cKT}�2h�ve����2��5,���1Oۜވ��4�5���"(� �ܰ`u�z'�'r_'�U��m_��?ƽ�) 3�n8A%����Wڪ��l/{������fM,=�q�?�c�tZ�R�{E��a���پ����]��[���#�6��n�i$jĺ�gИ������D��~:��I�����Z�6�5�E����?���K:��������Hw}D�q��hˍ߀]L.X��[nHr���@<ߎ�P�`q�A����D
�7)����g	P�/	����Olk�G�����h��ks�c`z�k�����F�0shlzs-���6*��7�o���6~<�q~s�b&*��2��`9�h�ޠfK�DPo�/t�ʒ��&t9~z�{��*�a� ����.f!����m;B7�|a���D��9%c������?�(��4�=o�8�I�q��b!�,S�����-�Ȝq�X=���P o�W)��ָkH[;&��kh��9\�9�ex*��RM`/�mK\r�Jobb*2:$���]!�l{~���,��049 �b�OB�0��!%�%���`����ۭ� ��U�v�	l�5�!>iڮ@l�w�n"��w���D��N�v�r�\��H�g�C��$�M�Ĥ<�ß��!�)�����.�ɋ��tX�Ƨ�;�[������L�O?��R E��>�!|)��X��;�Em�B�]�� �[�^���
'}
	�����ʛ��ގ�$e���|c���	��b���N�,	@>�mKn��("T��#B�Ccq��{�7	B^1^��ǲW�̖G�u�_��)�4�Z��i	ZP���f���I�	���szb��,�����t�ze�w�唦�^�d�J��AR��WuB���CLj:t�iS��J����G�7��*��4+^����%H���؂szByճ	����=_REfr���7Y���t�wa]��1&C�]P;��Ȕss�|���e�/�%��e�k�F��u�8�4¥}�����
�ipY:@/���Oꂀ�����Uճ��CdUO*��DV*�O!oa�,����~�ߜX_a�-�$�1}��-�<���<�Ad��}��������
�9��TATU��y��W�X�1�gA>�G��c�R�[���)b�nG�杊D"'�F%�V���	��+�8��be�H��٪�D(�(�t~��u�?�Q(���U�����Rf�$�,CC������[�Z��Q�"���gnP�r�j�ϕq�A�H$d����.5N���`!���b��Z�Y����9�O��x��+�}��U< ��U  7�w6��[�$�[�����סg$s#Bk5ݓ������A��S�l|3ȏ�%o����#�|���	B�P��B	jK��B{9�]q��1ZjC����EUɽ��.�^��z���El�;*C)C��%�uO[�4�A��Яx\<ɫ�ϕ׿}�ʃ/k/pa�[n9:��@򛽥?���@d�+�Ȭ�(�Ud8�!ݜ��!%�먕'9C0%|NI��h0>sH�qXI��q ,���)�ū�����_��!�̘Kfq��k�2�7�CD�Ë����'�N��]/��no=�,"��}�Ζ��lR_�.}�n�N8�C�F2;�*]w"!�Ix�r�I��o��Yݓ�բF���*�-��Nu�c)�4;IK��)S[<�A
&iT�Yh�%�ʱ�Ʋ]�ߡO�ʘ`��N#�T�s-��Zz�D{ϯ�1j�>��k�C��j"�� �A�ʪ�pڜ薊D�F?�_F~U-�?颣�������y����)K)�������� ��nB���`(Z(,$e)��2�K����7�8!ˬ����i��V���K�Ѭ���}LD�64�C���BD��ߡ_C9�#���.k�+	\oqm>(6󦊥b��S꣗��eD�(�q�}k�!|��L�z88-d�M�EK�����w����W��\0���-���-~ր��ծFy�0j�zh�)�q�8Q|)e �+�dJ7A�vH��{{�|?[c��#���P4�"�b1��'����P�,v�+�����}O>c@	}���={�e.V��Ra�\Re�3��{�
,���`ɀ[J���8�U�7�X�Q5�0n���GD6�G2���J�.
#8���#����ǥ�F����N����B�2���<.��&୽"���a}pq�l91hB�Ǹh��]UAc��hOMH2$��Ϋim�h�s��1W"I^0�4��u�l�6��T0���v��e�6��C��r!z�_$��?/ec�S������p弚�oh��5���1���&0�v������g��0�D���JJ5��M"ZX�9�m�;S�t�7;A��WG}�����M-zd�fj#]��M��5�b^��S���ݮn5�n]���	��<�KT�fk=���s�)���*'�H";��< e�=G��*���a�fdŋ�ה� Ye��fQix,��mG�����Zw�D���4?��<o�Kx�o����m��8Z��W��I�SSq�'�﹧��Ҽ���������>=~�qfp�Z$���_�4K%��M;�*&;����ƥ���aQ�n-8:����X@}��\ 9���7S瘖O�	��h:i{��i]�	e&��E�ߚ�E�j��mL�O2h��]�ym��Y�c����/�� �nH�;CFkJ��<$_z��h�\�>m^A>��G��$=��|���F�n�e����'���m3���K��@O7~���W�OBC{N5X����8���������K?��jh<%�F���CU�'�_�aOzȺ�#����ؿ\��o��e���:���n��ޥ`��a�'Ff��6���RB�xig㡒�Y�uP����UMǪ�F~�7�II�%�*�@��E��k�Lb�(�oj��Q�G�Si������!X���f��U���$w�Ҙ���K1���x^=��nEl_z��������
x�uMy����]9���C��(��A0vY+���-9A�I���_�n��h9A��ϭ� �Ίp���B�?s����9�۞oT��(�j���.'S�}d���Q���3�ӷW����0ʷ?�������7N�P�x-�߭^m#cJ�SG�ѯ5j˼wՀ���~����P�4�Óh�hlA��B���n^!�j?S*6�����m�<��a�ԏ���k
�4V�����>U��)�5x�L�9����3P-���r1 D:�sy�[bPZoM`G���  �YX���әX��w$V��#�,iz#�}v45����[�5}�rJ��X�D�E��XB����ʎ���ubtuE�8��	.I?��_����\mq:����8x��)��lK5E"|�%���ޑ��U��sZ��#`p���;�T� P��L0"%��iv{re�w�ϫ�ۃ���(�",�;S��B�P����zxl��M��+��p�|��(�����o�h���p=^L|nx�]��;�iA]�BO+cjL��:��x�{�~�� ��m��V�~P��/����g�I2��݇)�N�-S�����D4�Q$��AyNy��e����=�1ϻ��ۭ�s�_`B��4���q�M*��`-o:�&ҳ�%�pPdJ[1�������mIg<ǌj�A��� R̲V�?�����H��lB�<������ȅ��v`���X�pB�J3<�폸EG'|%	��27$KXܲ):��[kC$E}&>qo�? <���;O쮗-#B�����q�2��E栋})�{����XEh����5�z5�4(&O���+,�E��v�H�'F�(ԇ�K<a������~b�>�̖�J��F���0�Z[h��������Г]8:0��"��M�p� ��H�Ao�\�Cw�T�,���+AX�~N"�jc@�9���z��x�͛������-e�o]���T�=�г�ԯ6�#;,5��Ѭ>��>��� T�X�'�kw�ӓ�6Z\�K2�a��ǯ.��5�6c���Z�.�0}5�yn湕	�_Rž��T<��+U���Ϲ*]�c�|I�3�P�̽�Xt9<T]��SL��`M�x��a( ����.�N;��!�+e�����,;x��^��@
��H���J�d��?v��r5�Š}���o�͐a%�yH��{���ٽ�T��빩�z�1��� ϊ2��\>��Cu5��;����A_jNt��*���Ʉ�vZ��UX���Ydm����� �'!j�l��:S��6�w*<�]s#����P��%i��X"���֝�6+�����PĿ���}�Ͷ]F�*��Hn����lP��E��%�
n���~V��l�H�T�̿%la��v�ǡ.�C�ћI�낢����b\��7.�q<
�}Gm��r;zk�}�������l�{|�4	�������^�9�Mg�`�'���Gj����d_��?��	s��������4ȡ��ك�4�Y����W�mj�"߀�-�/oܙ�AG�	�_@���]���a󰼙�,��|W���������x��|>n��:�uc�ȸ�eǆ!� |0�k������.p?�w(�����a��6�vR(�+��c�;�2��-�܅��V*�0�n9Sd>�.y�/Ny,eՇ���T:�]��q���L��6ÿS+�1Y�$H��g�FyѰ���ghQA�V�a��������ԭ�$�G��#�s�K����x�?�); I���pF�
Ľ���6�t���7`+U�?2�!��ݨ���c �sn������CT�ۼ���3�/^uطEKs�,�� �Z��,@ӿ�)�H1��.2���moo�|T�<�7���s�����@'�D�Ϙ�b�*?���,:!Zm�L26��SB0M��91�jB��N�u�������.�?z�=w�cDfDZ^�̈́���1_DU�\�����)�˨P�I��H~���S�!�5]/"���`��2�m=n< ����!�c>lb�be��~~3`��x��{0�j8�}����5N����0�k5�t����8�|]O���������qv�-�H1�}�/0��WJ��:�4j������Nt�5 ��y]ѵ��s,Mŗ��QPB$��Q��8�s����(��Ϯsmt�b�i}�i�tb6�gI�b��ƢȘNY:SBj�AJ�k�D�ПO����ܙ�m��I��O�qE�"�4��Y�Z�5
?�mI���Hw)�@������d������]�\��J��{����w �)6�l�8�#�����Kځ�6;��d/Vg=J��������Ǉ>����H;��bAoj�.�؅6DE�F&MA�jW!�E�dt6,B���w�L��I|.Uwӹ�b6���Lo��h|�������=r쩕����������w͝/�Ts6�*��(7�K���i�hPJ�O&Cz�q�����m6bw��������5[�3�Tat;^���z� ��;9�q���Ӱ@3.�d�a!Hgk���,"�{��ר��L���؝S���7ã6��Xi4@r7&���P����I:���E��XWh�8�Q���%Ɣ��MP^�l[@�n��",j�a�'av�<{��@�*�{�CCSG�0��;�=�����Uldh��&��D�x�1�����H4���č3��k+���cI�O�D+������I%�*�VCݨX�sȌ�� �c�h�h�Mv� Zx���e8A�8=�+�"��.s�J�eSP�}�-bSc-F D�.&���1#�{j߻���5�?��멓�,p�eG�=�}����MoU��G,m�� z��d�uf'�q2�؁#��N��ѺUo�����M��L!�y���18�۫nzv�k�Qe�s���w�\;7a&�$ʼ�᪱+2%׉`�P���/g93ş�)#;�o� 񟜵�@��ަ�X��]`& �y�i���=|�+�n*�W�y����Ĵ(i ����+`<}JT`��s���%	��D�dz߀�PS:�ұz�Ri���@v��{	�-�9Y�T���!S��SOw_��B�0l�H���EJ����۷R`h�$��p_�4����3�Ά#Z羣 Do��qR�2�$X(������$�q&a��Mo�˽n�-��,�E��ڤ��ԇilq�d{`~
h7���Cnj����!��5�>�}��S�X4���{��1��A��gT���������o�����}d=����7�)/O��2�'̳��	lP
��9QYy6����,���N���g�x�x�A7�����n&z�Ba"J3!WL��u��v��4��4�T�����r��]�����SOo������ں�}���|���A��_/�z��cqwk�̈́�嶵Zs�-��צ�k�3,�P��z+���4K7�O��ȋ�	AR���UA�Iw��Ϻ_�����g��`ꖧ�����P��D��.^t���]���B�;�Z��a��C�gi�s*��$8@�k ԇ�O%��tW�	�kX|zƃ��jy_�5���U�Z��%�&�|�ŶaLT]&-�v�J����:͂����,���Q�L��� ��N��V.����f�qu�g���]q�1�*&�6`�;o�gv^�\q���X�'+|e��bA*V���7I�*v�赕 ��P��HSy�tJm$2 [�;��)@�D�z�׭S U���$11�4�)��T:i}`�����b\�B�B���jl̄���'@�@-���MsbS���gJq�lok+.%]�g���9��-+���.��Q,i�ڏq�K�Z
�{roo��f�}-�Jm$�%5h�*�����������Wnv�K�>0���.�d�W ����<]�����]i"���'�r ����!
���Nz�#��%�HXu�X�W���)�e����+֌�����@�R�6B-AؽN�g��Z�[�*-K�R�@�ǎ�	V�e�'K;����X���Q��y�H��c1-Rp��q��S�Ƨ��P�sҗ�k���g.I��z@���^���d�'5X��Ƒ�aR|��#�B1����o��?��M�]��3K�Ȉ��klE�oq&󑾼;D˞�4m>vt-e��a~����0
�}����s��)�����09���������������ܸ����R0m1���>(a��-X���_&Q����V��3bl�lȆ����̀D��[*W/��t�&C݈��x HQ���V=��8I�י�|��P�7'�������_�L����z?�䍹ُ�wwn^���t����Ѫ;��|U.L ������?��$��sє%��R���[�q�;9H�ߠ��&�xՍ�>������=�Nއ9�ME�b	���w){?��E�|��%s�Γ[�76�$�C�(��Y�U)��p�c���,bY-v�cc\�~lf�l�>we���%�#��

�9�� ��Q�f$df�l�ı)��b/��(�}��H�������(����T����;��͂H ��h�hB7�c+'�W���i�l��(�7�%�o-�BFZ0�Nݪ��Y�- N �w�Vs_������*�(P�h��)	��͆��a٤�T�4[=�������[��70.�!�U��Hפ1!�	����;����ҒV�d��?�����������J��k#ܯ���:L���.0�8gA	u�Kv�YR����t�_��+c�L�J���Ջ.h���#�Zt�c� XzµU�<50��ڗ_tcX-|�{�����1@�F����%�wF�d�F�D����$}�9o���S�����2�D����/�ޢ���d��9�ӹ�	Ư~̉�ȳL^{صK00t�^@�>RCMǢ�H�f#V��B��(J�	����z_����yr�NiiQ��*G���Lۄ��;�wk�k��rܖ��Yt��γ���W%Y	�Q��.G���ƽ���ό��b���e˻TraF���yQZ�.�'�����:L΅O�����aaLq?O�ݳ��-�whb���Y�K�[A�
n}}�����9�������ql�uee���m���-z!��lB� �g�O�I�q#�Kl@�0�f��=��A��P��b����C�4p��n�S�>�a�]��i`b-�"�(T�Ν��/&_94���<��+?��7���G/�/^�/�����;�??3�D_Ck��vc�F���c��iꍡ{�j��ː�N�K&���!)+�Nj1��C�D =��?��Ϻ��:��� 8LU7�E�&��w�z�}��ay{�s�ퟞ�o��WMN���hE����agҏ ���1"�O�E��.F��������E��W�r�LƁ?m��bT-@�Q�K;_�Y�����$lE���j�X��j�h�ٜ��4�@�ҭ�U��i�7J��9ڝz��Nl�XT&��Sga�4��TB�B��"�@ áx7�R4��A���!e��6���˓��nW�����(����EN�-�&�T<|�uױ)�f.��Y|B��F�I��,U34�yVpo��ä�����3��"���~W�c�\��5ʘ���_�u�)L���+ 8
�#-!� ��������v\�
�QpzvT��r�]��u�`���"� U������Л�;�6���C�����%��9s��>��MO}���y�R�r�&�9
V
��f};if�M�v�Rp�d�^C�W�jA�:=���cbtZ}�/������"�T����0���B���W�?�f�`��L���K�R�@�6q<3_]�{�uٙn_�.��Ƒ� i�(�b:u�X�	� � ������:�]vo�2��1b�޵�o��3y�/wv<Ţ����K�BgO��x�H��rڤ*��TA=�Q�}^��ʸ��n�h�T��@T�6R����=�S����m郊=�cS�OuF��*@�:���.�.��o?��C<���>��܏>����ڼ�?��`ss����3��^�����.R�ˀ�z�
�"otM���e�x�x�AӎV�M6w��I��r���Z�-�m�-F"e9r?Z����@���Ǟ����;vak�������Z㩡>*�p,ݦ,������G*X0re��ۂ	(k�I�Tj� �SG}� Up�N�0����/ν�PwjUXDV�A,�����o����Q֏#v�M����_�x6�9
�$��34<�'�D�@D�Qik��c�=v��n��m�m��a ��V��
Q��C�Wv+�J�!�d�S���dI���hU���!�J-b�@n�bETu&&D�S_j���&�xx�?͂Z��0ڡ�&��wy���b�D��ĺ[_^q;�>��(��c@�.���U�$ �s��?-MJ�^mQM���q�$ڟ7��/H�� �e��m�5Uɨ��-Y�g_�,�&UԨ�X,��z��
.�6"�n%{��\����)5��l1!ӟ��'T�b��PKkKbl���JK����W�L);�S"e�`��NJ,8X�Jp��A�1)�4�JܭA1��j ���>O�A}��3wI�m�6�⹪�-O�:��_�u�qz��r:��_��!�����И)m�F�[%���r,�b�Zbmd����`�i��N�X�������ӳ��sߘ��k�,�AM� 	��uKȽ�Ƴ��6
�u�=���AI�ђ����4xK#ڰ���?~��4�c]l�����uѹc��+�<��}>l�������f���>�Cj��5^K�Fz���h��a�W��% �y�\���x�K�S��"�[`4a�������*Ȳx���cpjb�>�3nz8��A��>�3dz����O�A��|�o����׮�M�)��YZ<�o�w6��+��/IM�/�rIw�8�1o�Z1ν-�Z;q�z�-|<�<� �[�r�|����o���C��D�D.)&�a�S	�0���#J���@����aő�s>~��ޫ�W�lsf�Xw}�+hG4�iI�')���X�d�' �`��4b��$�(kTG`x����<r�}���MX*ʣ�$<n����q�U���z�Z9�����La����g���+P�(D� �4�x�	�4��ҏ  M��N�͢]C����fUR暋���4i��g)t>I���[۸ee�:�,�WJjw��,��N:z�f�z��Z��^M��tZZZ���U�eXx��:Ux���=7�����iI��wI��;tR_sS㓮04�2��l��?��YZY����c�Rc��t��%b�7�L�0X)�B.�gƒ�����(��t�*Y�t�J�UQ+�lO�1O^Yz���9�h-"��8�L��H�B��ݤ�tQ�y�4�e2h�H���b�x1C�E�c]����Zd��B̔�������(SF,_a'��{�Q ѱ���@^��mV?��4M� ��⣅0��H5��XT������|�8�ri@�o~��j˽z�[�בRz
Lei6�X�k~ڒ�F�����-�cB��^�l������S��yL����h�cΛ\�=Ǆ�f���X��*+�B̭4�b�|ߎ�}bÀ�67^�ݭ.���=`��� t�R�H�V�:�	L�!��v�R_�c�x�X>��t!�,Ml�LN�)���l_J̫DͲz3��V��
��[QƘ|�'�,Ib��Q��v��X�(n-)��pc��L^#��Eq�g��0�>���N�v���]Z��m����`�'1A��FA�����|�x�r�?`#W��s�?F�N��,��sD}��Mv�1�Yq��a��K*��o ۋ�m�j�~RP���A�71E	j#�ͬ�	S����0	jC^�Yy���牁޷�N�|gf�a�)��<�gN�9��X>G�Z[=3#y�P(kW����t�0RU)HV�vM�*��r��JS�����vgN̸��玺}83�&�4��4��º�޼�ބ�u�27�9��(�򨍂K�u�Դ�`fq���ɪ%���y�^���&�7��J��ľ�}�ɗ]��Rx/)���A
���0a�X[�����j���XH����~}�J����ֺgq`�d��K�fuu���5=�5J�|oP�����A����f�4�<�K骋����fex`�-���[wn;��4'A��g�����`E�U���XĮ�ҭ/-���E[�7W�������琜�m�dN�O��GN�DNZ����U hiI-rf��9�nL>R�{e���޳�$҄�x`V�K�v]O�e1�$PB	0`BM[aQБ�,Q�)�\��k�E��H��yҸLw8�Rk���9�������:�!�b�q������Z�f1AUf��� ,��]��8lݑ#G�eڀ����b��ǿ��{��Q�����;����@	��=�b�m���(7���dtYA\_��>-'�VW�cL�`U�Pݳ8���`��T��*	}�dШw�+#�Ux���u�3ࢧ2Y�Uk���1�ԓ1�5��k݅JA���n)�%�����3\�#t�$��f�����t�Læ�1����T��1"	���B 	�Y����^t�>J���h�+h�L#�V��T���r�c�Y���V�jT>=��z��
��hSF����:��NQ����=~�{��n$�}`��d�j)�J��&����u�w����o���3���em�u#i �.;��܎�j�����F%���9�Ì�mZ#ɦa	�-={H��P�w�*��Kz��U��l$��	I���}�=�<��4�h;�C	��Ρ��ʡ��o�<~x�S����l������:���֑���n��ѡ"�B8Y����Ud�GY;�?~"1=ݼ�[�7Pk����� �n��	M�2*�a�[_^w����z�5���W�n���������Pgl�a�5R�w}T_��>����D�8*�%�VM�ڽ�k�-
Z��)GU�-�ώ	z,�;��H�Gԇ�t/L�*��L�߸�X�TW���!*�fX�}�w	K��{�iJ�bQ�8M�[[;6��TQ��~��̎L�8��?+ 1㈸)�.��r�K�w\��!	n|�N� ��~�-��'��0�9i�v e�+���b�hC��>��� ��hGN����N�䲤;,��<)(���_kfp�ɼX�3�fT���a�� /�/�s��F���s�M�wQG�k��W�I�$��,N+�	Z�vA��Ƀv��+S�%�F�	;(�"bM�&&����7���e��^���Ձ�~�;���f�4j��8�y���^�9���xM�އ���X,՗��{�a��˰b�G� �Q�6o�M���f�Dѕ-؅�{�f��\�?��o��o.�]�P9�o����t}�6�k��xd�`�&�z�K���P�2|���?�u���ҁ)�'��Y�/uJ�EiH1KJ�J'c)y� �۾����Ų��ȧ����R�Ļ�%�.�X0����^����\��n�0�|Y��_#[V_)Өx d&������*Em.���C���ydl�i-t`:��!�E������9�~o-��؛6�{0�w`���m$���W�<Wm5��%�����3���[95M�]�������А�E=�R*f@���f��3�m����/L�Rc�u~�C��Cu�y���\n���q�\����3��"h� ��uX�;�;��u��z�V�x�x�AP�S���;�,�i�>���ʶ3R�&��8���Ho��{k������������Ã��[��#�=����l��Mǹ�b'hMQfOJ��A�M6ݙC��̶a��r���
�+���wiz��; �ew��� +v]Z�������Z�0���ȩ*��
KP�R"�Z�����	���O��b�"�����B[�2H���l5S����
,��+�
���2�.]����&~3��"�I*C;�4�x1u��xk��J��o&���ص�A�3���.���u@�4LV��-�:��DݣtW��X��
:�e����;v����h��$`���1�!�Q����#����
�<�����:� Ny��2�ۃ��<�н�0��D-//[uN�K%����A����w�_��O���E�'�r��#�^&�V��!�{�%F'e#_٦��ZI(��r���2��Z���?���0a1�88�mq]��9%�`��n�i\�U �9�J��k�[Ȅ�%�$��B��h�o*�sea���Q��"�V��z��U�R��aIR7�����R���l�mn�;�)ֲ!��3H�V]k֎���>��k����ւ�TF�1@��-�V�ñ���D�qz���>f��P���Q�����ʐc�D�*M��^W��&$��d�{���|��@,�{Ü��{8�t��|�J̵����+0�	~�{��5�Y�W��tN�u�v�c���2m��-�ϵ^jJ	z�:֫j�ڀH��HR�Tal�X������6�{�j�l ʤ[Ġ��1�gT�]�^���V8Ί�ڔ�<��Z���5mނ�qOH����x�*G�d<��{����"~TA� 1e��R��s���<�sB(�+��`2�<*q#\�� sW���M*�z�r�)� \{���zص��~:��'��C�H	�U;�T�6����I���o�&-Q��|e���������M���1|�O��3���ol�l~���<�GO�.�����n��ւ	�Nb��~ũ������I��gNc_d��Ţ͍�����\�x&e��]��8hSF�Ǆ�RDj��^6eL���|3,�t:1J���x:�K5��d5{;}�ID�;̏�=��*;� *Wg��3����-w��7{�&�U[njߤ;��i7��܇7�U�|4��j��b�X�-߸i���R*������ Ppg��m��s�}��C16��ݭ�u�����v�B��UB=����F������L�s&u��=�QPUY�tUة f����ʩ)�(�4�.����cY�.�(Uv{��0#�]�� ��4@�u@�zyY/ړL����[��%U�6c�������)� a- �ˌ#�x-..�5R��^�6��rE ���t}���0h�(tF�����DՌ���KK_����hs��<״���~J'��YbS�����KћL~Sr;���p9ow�$H��D��.���2n6�N��cv�3=��Wj"�?~��m>����?����o������A��IY"(ĸeM��v�6d�q*����*�-(�d$fP���D �Mh*�x8`m��@6�mQ7�{@e�A�J�Go)��sls��^�g�?�K����w���A1����1m�1V�)ɻJ�`O�a�U���XY}�A.�丬c�Y�*f7b��tFO�g����@��D ��� cw�?�&�G����b� ��Jȥ�y���dU�S��&T��(���yqMu� �m۰�T�ж-fW��y�Ҏ�6�|Ǫ�Ab�p�b�5=:��'�����]`��N�?D*����x������8���[fL&ؐ�:��u䜷T�g�Ě�|����'�����j�kG��
5b"�XϷ�0�X;1-���qs��i���y4o͌�*k�������l��B��J>_��]w�v�;�ɦ	�5)'��.�&�-��C�sϿ@�g��h�l�&\݈K+k���p{��v���E��hRz���"G�lx����8��y�'*��r��
����˃���k<mJ�DT����x�2�Su��E�W��i�I
�Ͳ#��}�^��wX�K� �6�z�Q����&4�_f�j�P!���8����'OZ����h�!/�n�4����8��~iR�]����r�.T�h}� ��-��sg?6/���}Υ{7�x1���>v=�7���4l����L܂%*��P��؄�]ق�(�҈�0)�R�+��LL�*��Ɲ�t@Ī.E��fV�5-,
n��;�>�2�3/���?|ȍ�c�������GcW���Z����{�*�A�m����C�Ȥ7���J�#�hqx?�%����~��!i��5�� �yR���ꈛ+Ɣ����g�iR�J�%1*��i��k ��_m<`�`�tݣ	�mE��&Usy�Z���=ģ��L.I*E�YL �K�o����\n����y�"�� ��@G�t"@�hsw�=�Hv��/�Ο����e�X@y�#Ǵ��
OC�-f��ՠ�cK"��V:���Z#,�tIC����{M{�C�a���m	<��D�H�IbaKsٳ�M#�P�,��}09������^��<fvN҄u��Zz�{73����6�#������`cgk)Ƴ ��$R��=d�@|f�]����ݾ�a�	҉&�9�4���P6�v9��ruXCJ�lӀ�-�3���N^��O��I�SV�͛-��q���B6/)���ᓃ���̟��ط�U�����q F�6sU�6�a���Qc�0�(p�yy����U��Z���#�P� r�t�h4y(]B��B��Q���KT��|xvcjddn��΃���c#��`�\(n�s^�r�<k�s��#�i� ���G��}	(����Z0��e����'L
�cW�ᙞ5�n�:��A�N�� �Z���TA&�U��Ywu��y�& ?���L΍,l��Zh_���b���m�4���0NP�n�r�n^��MRe5����Q�KC��ַJ���2bf�vJ�S,�ڱF�8�~��`i~��^��=l�c0#��m�o/X�����Ыj�}x�+�6]�x��gFO¾���`b��gM���82�RG���[�n�����wp�E�V7��<ǭ��%αH:��g�v��'���kn�j�i6�9����, ��/-|Sv���6�y��G w������)�)�� �䤥�0rZ��,&�����g��G�̵JH�><���v׶ݝ�;����Zk�.�L-�Yw`�Ǫ�1�᫘�#�N� ���yw�8��޻���p'�uüW���F�%ؘ("�dM�-�3Rq�����j�
��"�!��3�r��⍬�DK����9'�!i�~ ��Q�ɺ����=ƚ��ԚD��o8{��ec4N %D�FR&� ���������6�w>����YW� �1�S���k)Z�4��8Q�(GkURZ�WKL��|՜U}I�c��w�x]�J(���WB�<�
	,	���z�I�xX��&b����灔Ϝ��Fac�/�a����B �����l�Fbp�gW3d�&F�૔Q龆�q7�x`������=�BńN<��K6	$`��
���Cn��g�t��CE��	,'&S0�g�������<_P�6TAg�������t3��'{��q��y�e	Q \@'���Kf-W@�)az��ET��t[�x�x�AN�=LD�~��M�Di"���<b�{&�4�{�>ߓie��8�|?�0����1���L�;�
T�����I���j�q��Z`$�ʈ]P	�(g��9@��.)&���^�L�0��<j��
Ti�7BZG���{� ���,*f�dS������;H555I���D(J�����;H����_~�e��U��z���ܩS��|Ϙέ)vU����>�2�숛�d�/���vY��%��H��sOMOa��Y�V�mӛ��9d��&����d��Y*���~�Q������۷a	�6	��c�臦 �2��,dm(�}�y��m�o�`��0%��Ԩ[�x�56Kn6F,�<��j��Q���Ӻa�DPi���yw�T_�pϝ}��I޿H�ha1��1e��{ ���J�k\s�8t�s���E��G)P�>���t�T�]|�R;�e���2�k��a7�������[wo��s'�ẜ�f���K�����)�kBŏ�_�6�7Iʋ+ @AQ4�����!ӫ���x�`��1|��#��k -�_�*K�a#I�d� (%�޻p�C�t�ҩM:xۂ##G�-؛�\����=e����7]��%1BR�*-k��}|�!Z�5�5Ij~P*H�ͦɱgI`��\�Fi5�����w��"]�keاԏZCt}~�G�������l�.����?�qb�@��e���9L ���X�<�2�;���⬋���n�ژZ��]$�I����w�{p����DJ�F��}��M�HQ��m��l���-�V5�U����^��\�i���f�/]��-m�=�4:EY�{�KU��i�MU���v��B�. z��z𱊧�0F�����P\8b�p�:݇z=~�����P�K�]���8
3�c��.��iA��������k`��)�0x���N0���yQ�VIA�����=���)����*:������;���C���B���;�<��2��X44KL���&�p�;@�)��fH9��9���N�L�^/1v����%���m��H�A������v�������D}�F��Ϻ����a5vGV�'�`��2��-� ��X-�#�V��۔̧��x�$�ffbj�mg6$��Gn�Z�Ϝ<�:��mX�=b2ˡ�t���c�z���eU��C3�����ʅKɞsX�&�?�ު:=j%���LML�W^�`���7�֥�nO��b`}�:�@� ��U4�=�~��ť[UX�ˈU�Z��c�]�4�nزhu��T���0[�MR)��O�c���֦5�]]N��vؼ�� �F�oH�,�g ]� f�8���hU���ɒ�:2}��r�67�G����+,�<%��bb�����`DN�jC�d/���gu�O��&���rW�OZ��0�-����Ѯ C_�����+W�9�<8a {�TeRB]�e沷@���5~�����G��H��N� Rw`z����^ ����uW�f�Ʈ��2�I�X��$�;1���is��K����� �IǤ���[-c���ZM�Ě�7I����X�� P���J�ɨ�(r�|�w,PUJH���b[���q/�$���=1
ּ}�ՙe��X�����,�4�SG��L��$�M8�تWW\�)6]G5���sT�1RR���[�bP�cWH�2'M�!I�Mw���ؕh�TuK�eR��d#����'��Ӝ��8��Ο���X&�k_���%����c[�~WC�E�E�Y�@��<��C㽻E�cL@���U>�� '{����~�%<|��75"��UEi���ļ!Y�E�C�Pk*���C��c�և�79]B1���}(�T`�ːZI�$&V�Դ~���ƪ�+�ϸ��_pZD�Gs��`!���굛����p��XT�;48���ݸ��L�tF��K��i�������Kp3��ٺD��;.MUB��C�*���Μ��*4��O�xa� ^?�.�{K�����W_}�H�/}�����M�*� �{8[ʮzRT�P�x��0���Q���i M�t�t-�Y�=X|�Q6~橧\�f�Ʀ��<�n�"RU� ���+��s�K����⊹E��ŏw��c�,����8MO5f�M�&Ww�(z}�|N*O�y��k��aw��U���[MB%�|v�n]�᲻^r�������XK��o�!��f'9�f�}�Rk�+�B��B�O:�2)LU�r��G/��ѡn����uJ���t(��J�Ro���J�~D��U3�TbBN���ԕVDp,O#V�^�� ��}@�t ;��R�]A�λo���3�yڝy�q�?�� yc~�m��-^�<��
��i���4 /�}�A��	Z���P9�5����V3��RZ\¿�(�tgZP��*bL�8v��0��B]��Z�:NiS���A��9T�t�;h����~��;�W�\�^ �u�0�R�\]L�0�Rb*�V�R�>e�bq����'�P�+�d�y�f ������@R�%���Ĳ�ٴ��������@�= .�Ǟ�����KKw�5��I�$�G���-Mwwr��y� O��%�zr7}��Lbd~�H �����k,�٪��m�,��H]2�ײ��Ry��v�9�&mƪU�W,�Ƽ9��)��S&=�,	��(U�}>�A�u�ڠ�S	$�oϰY�)��R�Y��Z�����}tij*7�v����[wfL1�ޮD����1gk^�ꜹq�ʆ�������?���ơ��1�I��p�dAϩ�c">Ɠ�rK�j|�T�%OM��C�?�,�Y&��Ivd9&�Q�<z��G��yv䴝�9lrh/?����_����8����KKn�����+0�eԹ�X���AT0��g/~�_~��-d$`�Zjr	�����Dƚ��r����\�r��շ�>{�=����_`���.���ʨ��$E*�e����o~q�M��>43�|�3��n�&|������hC�#-܉�����U݅6h�Et�#O�qKsn�� d����л��g��z�r㽳
���f��!Ť��L���a�{�T���q�ss���g"��r�5"�}［}�>9�n`j�<~�J���w߄��֣ �R�M �4�F�6oܢt~ü�n]��}�y�{�J���z������"��_�-i����Νٛ��7�vEؾڝWǏG,���i*�f\����p���Tr�ϴ/�X只(����H?��@��nU,i�:�D�*�|�	��#��%uɽ��{�C����;v섛�9E�n�� �*�"F=�H�Ŷ��p�u��6��eN�$ GQ*��h�
&A��"�Ey/�^�f�Y0U�f=x�@���%����y����o7�\6p0<<@��Xt�$������~�}p�}'\-F�W{r���7l=�Z�]�������*L�~���Z���C�J���L��E�-K��XQ�}7u���^P�%FP%v�������?����݃����G+���a�ed�)Q��_UU��B�y꘵ȋb��D�TmV�\u�����v�-�K�w��k�bj�VߠoX���"������K. ���,��Q�A������Z��9�����'��#�����{���"�	gڿ���~�As��
	�5���g�z3��>a��h�x�x�AP:��D#��[����g1?�̾ƌ�Dm�?���c=���g��N��!=�~6w��0
� �]�a��i�-�IkTI?(ğy&�i�����)O��2/�LQ;�+�/��/�5��F���D�~O��3Y�Ƒj��E�C��T&��o������@?iRv�-�z���j8T!�g�:T*�V��n���uR�T�9_������R�U+�5��ƧM�0�jr��d>(6I-,�樔Z^t� "��nSY$�p���#2�F'&�����D��D+3¹�U�JI���nGb�wuAp���i� �SA��~�`q�[���!@��J)x�$i=Z�p�#|f�&*zj��n���[�_���:�&�>ۡt~�0�I�D�{�eݡ)<�hH�q{ɍ��a�����<b�u>/�8��*�nR�6�>}��"׾O=�X�O:��h��ֶ(ק<W-�
��EI�vI�1a�������Ô��KK+V�6� {�$3(�F3Ō�~CCL���=r�.���U��+� �^pO�~����p�I�mo��/��-ز�LT(Ɠz��4�R�Xl)�T/�4rOEi�H��Χ ��������O����|XWq@�����0Z}�.���<������r-X�Ql	~����v�`F	����~_�>��/���Zl�w����g�Ll;z����	��(�c���W����|�Y�/MX���rF�Hs䁊�9�t�\Q�$��o�j1��F���.Grwj�f_�k�<�AmKt2�l_#JGNlD�i��b^�#k�(@&(J4�1�K꫍�;,t
ᯎA)�2)j�!4���F� &@ٿ��S�:y)m'@��V�Ƅ<�`�dNP&�F�pz����-E�2O@R�����?��ݟ��Rq��6�v#��g>uJ��ұ�d�VS"|<�<� �M�H�N��m�n�a��~�l��E�Bڍ%�6H\,A(�9�:�,���Zl?���I>N7J�/�]#�������Q������ӧ��z���Zy,��`г�]�t�}�O�'K���0��qc29I� F�9���/��
�S�N�q	ć���dh�&A���������֘S�:�K14<�p��J۽����W�i���0O?��J��G�D��cqʛ�[�wH>17���i����Ѽ�H]�Bڊ����d -�4�������lZϬ����Gƕ%�>�]�r�42��Rm&�t���;�n��I��C�}�%Z$�������q�|X-L�Zl쬸�oߴV$�2�9uܝx�q��]��
�g# ��{
�S�]ZB�:�1"b䅳��܇LؽK�T}#�<�a�vC��GF�8�|�6��Y	�p�^�N�ںy�b X�ľ�Iup��[t�,�nr�4ڤG�*�I��n�J\��G���,PUw�._t�&@?�.}�V�̿JJP�3�QPE�d
9�C��?Ȱ�C�B��ء����}�]��Ywq���>�溺�����]�`2@�*�Fq@hC�h�����Y���?5��;��}Un�w��Y�Ӱ�W��ٔSsT���r#��|���J�XO0����U��l����k��Ywf�����:�����9��@^���x�*�N������k���UIzt���yY�Y�����on{bH�_�*-1!&R�~^h�fC'+���YU���`�2��co�k���X���r��tA��P�:(�$����3��n�GJ��?���F�cE��	H&m�$�ZA�E겊3x�L�����ީ)��_.>i0L�-�CUyId%�R�6�H�,FH@�4�*-a���g�x-��8�B�S�w���?W�Z�����Տ���ړ������Aإi�3/Ț"�E�Xwm^�1�bT�� �o�O��5J&z�k7W��x�N�I崕��0Q��	!�g��c��n_ڇ�os~������&Ŋَk�/�?[�z���XV�� )�CFܯ}�i7(ֆ	$롶�o�#��+�e�?�"�� �@N�	��x9A�G�]��Ճ0D3 �(Q��Xw��n�0�;�+Q�%B��Ha�LO��r{��H�n�����/�#y��L����߁�E;Mi�l4q21�`��,�!U4��_�k�B�*�9��z�S�|��c��6	g�6c����B-�@��7�H���>�/+�`R��Q�4^=ۀ��_�t������M���:� {��» �B3T�������ހ�!���kp���y�X���6̃D�	�U�(���?6�
������$���.e��گܦ���b��h����O�S�H!�7mS߀\���c/>oZ	�т'�z-ieZ �>O[ ���$�)J���u�ݏ��E,���M��!t��R�ϝwح�a�뮼�T��α"U��S��v�,��X�`�2�?�;�{�� <�z��ܩ�ܛ���
�,�G��{������G9��[�u�#D!5��(��-�w�Y`��l^]�=4`�{#�v�H��Z���Bm�j��L�hy=Mg9�`FW`��?�%F�`|�a�u�[�A��?�z`Ӓ�c�Z��Ƀ��O~�U���.n���lTT�eU"g���WK,�R@&2�1��`�e��{+��UV��~�E�g��o�4��ĴB�h𜸴JJ��;���᫧�P��􀜷>KvҎ�3��x��I�n�z���&U�u���a�����L6 R]��9�������
��b@�,�����2�#��s�l��*]6 v�ť�xaD�����2k �
�Y�Z�IQ�Y;����L�n�}WU��0q>֖��O�� �^v�~羟����7_5;6�	6xq�Db�d�8�� ��\I����>pj�XR�����톧������Ve�^�+�-���1��jw?��}�ѩo'"��|M~��1A	�H�$ 4�$G/�~3���[��rj]��?T��Z:]�"h#̡]3�9>�f�EX�HQ-7(R�I/Z��S㔛� D�YAs��-����$�N�<_����iM�-D��w5u@N�4�Dk��[o�?��h�ÿ�[��^��g͔n��\�qM��fɪ���.�����It�Îqym�T_�=���*<w��,�c�ܣ���Z�`|������JF���P
I��i�#�g����w���͏?���mZ���M��T~���F�T�������)Q�q"��,��9�%G������s��6H)]����;X�ltz?i,ZP�������T��8x����I�&U�2�w^��{.�bv���枫�lU�$����Q��Ao����zt��y�����%�U��(�B�m���^��|�E��&������>�0`u� ��aI�����������s�	����}����ǰ�#ց>[�?4�]s�b b��2ڮᾂ�������_w���㏝q� *�E�	��2m"f�|qI��V����VK3�d����Y夜���XlW��D��J��81>��3)S'��r����[[r�z;��0���Z��7�&Lؙ3�����gݿ���u����fE�r��>B�+��E׃
�\�'�������7:���Ș
��@#!����":S�+c��_]�%sF�/���,�F�>�%ƮE�,2�n1�4��<x�txVZ./#��4z�#0a�U�5�T��}����*�s5@�1��ps�05�%�7�mIS�����=�f�_�L�{4׃�Y��������P�.� �#���j�=Fj����@9�pr����8��������DT$����?�����M�b�Xe��*Y �F�*�a�jRǍz�O�`·�	x�A�X���b� ����(mw��3U��ͫ2�v[1������n1y��ke��3y��,n��hr�|��~�Z��+��?Ja�:=,w�qR6,��(����~�ޭ�/���V��oI{�	b�#�OhhR�I��bWn)
���4�&��T!x,�[��b�m9�,���+ ���C�ҫ����$���_u/|�Y��%�ȺJ��MUc֑��*K��e�����^ť�#�cK��C�zVN֘���/Q)D�F��p�0	,\b���e����*T~��/�n~�ł:E�L��3����aZ �ĥ�co�1X�ս�{���z@ x��� �u��*���<mz��!%06��v��K[�WfM��� DS��[���K���9��j��=�1R��c[:t��B(-,��-\�b��
��S��_-OdP$�փW�R��)��""�2�J@v�/\t}�M _�)�N�CZ�2is���Iq�#Lȫ��?�QJ��nK��j� æ�'C�^<[ġ �J�Wy(�d^��GN?��ɺW_{�}��� �g�u�&��0�Z[���#���G��� >��:�ے+�	�����>3�L/Wo�j���C��q���F2��\�]D��,�q�%řU�L^S�W��4I�@�AZ�i���%w}���HU��P��9wSd�jJ-#�d�����̋HKﱣ㗖Ơ���<K���tZ�.������������������_xpe%ņj,��#k� 5d���G|Y3X��y=��a����y�<π�>����O�鵘c���G(T)}�7g�O�&���s%�Q�9��[�X5�����V��(��(��M�|��
���9�_PTo�~��R9f)A����4V��}T�=��YL��ʰn�tk��ȹ��̲������ez�A�9I$�U��|#I�7h2kr�VIm�I��ڣwF�y�[��x���kt�����_*&2�����k�/�mK���j������z陧�����r)z}EXP��d�8%�[�fᛷ�����A��(���Y�32HDo38(��IѢ@�&��Q�M�ڽ�o����� JB�K5�*KƦ��FhQ1�.�fR�A������?�Q��E�8k�XQ{$M�9��ի4!�k���j�;n��l�ĭm��a�<��;n���'`}�������ԝ~�q�~ȭ����S ����7a�n]��nP�$��#�=��� ڞ+W�"6�O5��	�_���//.�3Zu;���W^�R�1S����Y����m�Rl��(,�4�?= �y�(���f��j�L���Y���{�
)�z�5ѯ��\�� u l��b�3.ѵ?V���H�0���"�+�D�t�a�҈��c��$?K*NME[�N���~���^��j�١L<õ�e<l "Kw��ƛ��l�3��	���_]��
!E�.�;���,�+h����n�� �R��\�<IϭS�O�c����^{ �����Y�_�uw����L$q�Fܾ�� �Uڒ8��z�I��Hq���g9<�iA��!a�f·�r��0�2�D�V�;yU /%�����V����Nsn�@H���,����}�}�o�o��1����ʑ[����ia���1_���+L�x
���WGY���:mY�L��SD���щU���e�L��@H(K�&�Ù���O��mP���|�<콼�ڋ�}KK��X���8Iu��&��T��
f�z��{���Z3~��Pgj�!�OG���$���+db���F��Rxm5}Uu�`���9�(����6>�˪�b�S*q<���N�[�~ h�з����J���`	t�� �?4gw�?��
��]��>�$�]����W�߽�ڠ�����6oӬ��`l6Z!�$����Ѓ ��m P�y���W��d_e��C�P�ڤ�w��e�S"�����|��)��'�����y�>�_D���+��Mz����N�v���P�(,B��M$#�c )i�n�^�����٣�a�&��h*T&&H�|�x��`�{ Q��=�M�k�|?��0�[���2W���O��J�=Z����6?���3��s�
�Y�,*�J%*�8����Z+���#�
C>N�5:��W }��l�`C���2g��1�3��͎q��V�>��s~|��~7zꐫ���If9�ac���/�X��*#�m l.����?��)��@$=�y��UՆ�$�Q`��5�QsWYHW�Wp�F�36��y��F:l��G�
��J�H�Ȍ�_��*��:��G B��đc�Egv5h��v�M���j2횻���4�����n�Ԥ��$r�"t��z�I*Ҥ/�F.&�,�&�(�+�y��v"g91mϽ�"n�����Xĩ<�A9m;`�
C}nbl� ��K�B�x�SZhi�E�q�Sݢ��H*��l���ش@�� }?��V5r�V{e]6 7=���~ޝ8��ཷܟ��G������N!^'�2�܃��q��_{�6��)=���y &���+� K���R;�]��)��^��p�?�p��i�}�rMS=�,��W-"����ݡɂ+�ʋnuc�}���+}]��W�ZlhV{�n�e��t?��t���w�c��}�"�Uc@)��V�J�=PL�@�F�U�*�W��4B2��6A� Z~=f�� k/�?���a�VgR�Gz�&�#0'�!	���ǂ,�V�c���d:���ڪ<���Z��(�H����J����_�V���ޤ��b���4�XU����uV�2x�h���
��N.��-��Eh͢��F�13�KK��*0�.{��9*H$�q2
(�c���G��?nR���Πb�������HP@"��.��D۴��B.�j7;���#�Ѓ �+(0;u��ڕ5��tct]Tm7��� �d�X��X���vo��~&��az�2������Ӽ@L
;���7���>͗/�%j_�����es�5���D�*J	��ͷ�-�;o��6�2��e*'cHڃȄ�Yk�EH���������YI��� HFf���3��@U�o;�a�"[�k`���Av�	�8W�w��]7L��L�$XV��aaJ��$�tt�~�C���FB�"J�h������_G��N>��4iR\W�\�����w�8�Z��ĢeìR>�c�h�B_�4;������}�p�"�caU$��,��8%�'����[����O!)�äѲAL�0='�h�
�P�1��3�ƕ #W���M��Q[����{��+���KNw�_D �I>��T���5�a<��O�t����K�7��-����,G�n�)RA���� 9*���	4WC�a�i�я'�(�yP�c��:F�+w0.�s��h����C��m�Mw�<A��SL��'��r�P��-藈�2���7�S�pL01g ��8��Ť\��= �2�Ǳ"q�Zo��ji��P_;y5��֍�o���R%��/|޽����L�S�*�H��u���0�UH,�U�e)\�U�n�R &�M���Hu�����L�t]۔��aʰ��u�_����|��o�ȊR��ޓn&�9�vqN��~�nv�/���,�[`���K�#��0� �����ӑ�����t1�HB��� �x�4�J���.�*�ׂ����`3�U\w����_��Tc<���eY�|ƻ�-���w��dFV�H1w����D�U$��T��34�>��O�h\�WE�\��﹞�Uo�ԢQ�}a�tn�舅�s�=�t�*?e��m�`V^Ch����x�
Vљ�b��ǁ���%�����,�l6֙Tn�Q���9��[��>��㘞����]�?�O�n��ma(� �����*IX$��ooD�����c����_Ta�@��&MM�I(,��g����D�E��W��Έb��#���f /<���>��"�3��ۼ����|�J��nCT����I�������t�EmC �~`mvH% �Ǥ. r��0��K�&"!/&�d�M�4�U�h���KN��2xѸF)�̦/n^ܚ�Y����&51��j�!�m��,�����ZKc�� �ߗ���&e#���GDz�~܊o߾e�eme���6�[M�PF`]_g��)�~��zFz]+O�W����U��qz����a�no�T ��c�t�7���ܒ�C��<��x?��4,R�t�0��M�4y�q����ФWR�����I�ȋ)K�j����!��߇�6�s���:USQ*�\�l�E�9N{�F�ucڷIz0�I_T��aW�<��⅊���>K���4��!,�o}�>)�	W/�`zf�� �~�c7{��-�9�E��k��i'I���H=��{9��yw٭�|��M�n��xI�ZZ\#\r3���)��QS�	u��V�<dZ�g\���; ���"`N�R�����Tо��e��R�Q�6-��;ڋ�^T����'��)���r�#���Ym�
�~���)V�[)7��,�����SbS�Oβ��T��i,"���c���Pʯtu+��~M�	i��%(��W�ZK�c�d((��~��i��o�}��[��X�\4�-�vFj1��U�H�찅K���x����\��q5�[�OZ����t::-ݪ2Sz�����
3�HK����bν��y(�Kϑ�ǎ�{�æG�����[1Q�N��`�偎��Tu���8���[`E���D���qo��*.6R��[���9xm�d�`ZBm�8& U�9	�>�DR�pFjP>�m���@5�{-ڠ  ��*�>{<'�\�6C��l&6I��"ϩ3�` �<@���ԧ�O���m���g��\�m�u�D��qcG)���/����ZZ�D-K�k%���o厬�f���i���
�1[��A�q�����{�YD��K|]��/ Z����_������I�(lr�,Ҫ~��K0  �+18*e�x�
�W��-D�T�0�!"�	�zwI���^��2@�W��I�VX+Rݻ���Gys�*�[��ҮR��1<`
to0������s�=rl��3����=Y�-i�\qR\�O)�}�զ�')��x`����"m$��6��ϗo�q�8(=~�atLv7�z�-]�,?��R9�p�&6ߩX��1J�pp�(��D��E[�%�������>�Y����c�J�X�*��9�oQ��bV*�]���ıP������]��E��Ћ� �g���ܭr�Q�Ι����9Be5��
��
,؍-62֚���;��ݸ���KEU*��q��;t����<>:c)7�;�)D�T�)]������62�s�^0�
�u��B�U�Z��oz��s��<E\z&�܁bƍ>q���gD9�u줯�S��gurߢ>�4^�9���sOp�C�<G�m�r�=>S��} ��YYt��3&�N T U2xܦ
�O�����/�g>����^v�Ϳ����|�W���`z�Mr��iȺ�U%}��(Š,���ԃ,bZ5��Q��Wa����e�!u��eP���gS�X	tDH���Bkt  \���t���)�K#[X�6����}	�Iý��%�V�21�ܸ�#,�f�Mw�v��1 �|❟�:kh�H]�	zR��E�9h��Z�(���T��{A)"Y/$��y	��U�ܲU��Ԛt;�q����d���7riF4nP9N4�M��yN�&���-Ыc˩�;����=Uw�T�i�%���#F��c�������
�s`��L4I�,d�c��Zbt Nf}h�t��T�K�x�wj�Q<�Lu�M���^����6����=�<��؆v�����Ͳ�qnݼ���#Ч=w���'F��ĮIC^�b�b�Y�n��۪c\���қ-���A�{�����Ѓ ���e�^J��|a�|y/���D�1U�����pc>Z =��t�p�n�e��Ƨ5f�)���|�/~ �giG�IC�u�����}���i�ȴE�3��/�����b62T$m�o]����Ź�i��Gis?Z���7�A�5v^F�k�'�Lλ�0@����u7�8O;�RJ�7n2���W���?�VB�IT,�:f���"L�ZMD�~��P t<��ch����'��
��k���<�V���E�}aw�i�c�.�� E�ٳ�I�_0WA��
���`���ˆs�?�&O�R鴼t6�(Sz�珲�Ϟ��nQu�J������Ec����z����	9HZn���K���-_u�M�W9R��֫�$d�Q�E��΢ c�g���A��m���/�������ƻ�q�@�J�o��=�E'S�B����ep�����<g�n�M* |Յ}�(��M�MX�e���G|�CL�-���"1jV�V�y+��[���͑��~�g]�F���_�w��{�ؾ���he�ܡ�q��{����j�:|ش_)t3M��eF)&A��`a�m�g�s�\�3j�ZȺ_����m��/��z���i�q��r*1~�=k�����\��:� �o��x�20� ���6ʤ@�q��PF��~������C\�Y���N�Q�k+��)8u��~�4Uθ�ʇ�W�dqoÖtHJ��f<��ܺ\��kL��je�B�C�,��Y���IPefˢ	�I�q29�Bo��9.U�ɃI�aF�e),���\�T�m���%J3�zM�WUi%�v��{��������0ɴ#��i���G�a�U#=4.#��,$:�ͺ�c��T.��6̀�1��2v]�z,
X�N�vu�2@�2n�k�LM4�-ҁ�`���*��5c��|4Y�|���xh�zt���-1-�o�l���`� ��m��|x�o)u�Ąo�qZ^� v����I��@Xn.�������z���O��-I����<r0*�d�CI�U��[n������B�?��w.����aiu���&_��eB�]���?]���\�v��f���uQ�܎{�טg���LO���ko�Xo��ꓔ�pU�HӇh��n�?*uN�D��!��Ӵ����/~�΄�b����)�� �Z��Z`̩G�/T���3OSU����^��zK,F%Rr�����l�(u�*$5=�1a@��-��XF+r`�(�i=n�w��A1�c��?���XD������oō��'�9y��W=�6i��+�\Sz@��<B�� }Ȉ��ɑC���ЋI��\O����7�r�Y8��n��>7�o��;�px�e��dI�䙨ӅAs�ނE�y���7���j������.��҇����Ӛc��L}<=������'���G�+hn���?Ʊ�"C�1W*%��7_%�*Q�8F��I�N��n�	t�E��8��1��bM ��u��y�ui��m��`�h����鮳�n�F$M��+ <@�o�]��S'����)��c�l�n3�����6=Y�Ta��aK�ʕ;���c}@_��lYy�J�q���k���B-Ɠ��K���[\�vg�]���( ]��tc��൫���S�X�B0������V,�R>�q��'Cܫ��b��$�PL��o��W`tz��b� nn�(�'5���:`�M�ڮl��Ȼ?s�8���.l>SbT>�7�ا�J��~z(˻G`G~=0 0Ko��%
J۽������ FUƦ��6b,���Tj*����೬���\y�X�zXk�*'x������V %�2s���{�x]TUr���רp)�#�b_�)�������Ҽ��0�J7��0`�R�(�"��6���ژ�����?mz�"�S�I�t�}������B&�J���Y@P��m�[�,�(�<"�C
��a��u��"���l�r�����#� ��R���?�)�fR�ҏ5�'�wt�%���7�#��Qi�c����?݃��"�Ѓ�z�^h��I��RTMA\U&�:����{�S)ʍ�Ll����N�O��n�(J�J�H��щWOg�I�yl���� U4P�eh���T -�	h��L%L>JE5D#�ݡt�F���)�/��A�A);Ŷh`Z���%c��B@�)}�4��1�}3,<�t�,�1r��oQ�v�5y�2_}�E�AK�PI�lo��P��܉Uv�����,�rq>J���:o4��c��M��.�֦�m��N�$z�I}���%ZS�QM���c�!�4er;׬�C���%,�|��� ���Ъę�8�QJ�o_���3��r�ֱ�u����u���~����BsҐ��S�t�*+�=�	�h�̓�h�ܼ�nSB��f���_��YPeD׸z�%�Hw�*�0�7Р���8��4�e��%��� �u�q�7�͸�C4z��s7\�����,(���t���\|昛p�`ƴ�䯟uM*qo�Q�?�T�-}@*�����	���]�a������W������a�Ň(�@����w��5�j�k%�@óM1@��;�ɑ�C4lL�ݻg߳R�n�56��d�N��%�f=��b�z��\��t[������e}ɴCr��4�	H���%��+�"�E��
������ϻ���_��{�����cU���*��m ^f���83�Dٶ�������i.��Zq⏭A�Y�~��H����2���HC��H#�����.	J���Qzۥ�4UEL]�v�y��awVr�n������iP�ۣ�����U�Y�����8W�Ԧ?�o������3�3j�,A�|��Ӄi�y�i��ȋ��(��3���IF���Pz'	�k��쉹Uce>H:7�]<��)m��=	�x��5A�ؤ��ā�*7��; ���8|����l$Sz/�l$�m��3SH�����2X�v��r=��
<I$=�R�����Q5=�6�ܧ%0��橝af�Ӊ�/��b�0��p/$�&��29��(�}�E?���]ڎ���	��΍%h��b~Ԙ���A���t���*���~�G��ܦj�����u�$��/q�f����dl�a�QC���/�\I��k-2()6��6�\���cY	_����C�؍��K�f������z��#5����A���}q�]�Býsu��j*�OdY�T`qD�Q%!����*?�J��u3H�_�����I@�H��A�L{���$�z�ĭ]�5���_��5��SIӔ���L�)�YI5����\D(;6{VU���,.��r��] ��;.�|=-��j�S�GOT!�>�)Rb�̥ �?Q��\��)�z*����{�������r��>�GJ�)�8�t��� G H}�mk4Ŝ E#M�R@�$\EkT�9ڄ�S��/~�:��Rrj�8����)%OQF>v� ���U�\!���߁�bq���/�{D6�1��dQ>LW�'�\���Q-CV`4� �+x��W߷�m5UϩCGка�4S��W�>N��v�W��}n6fa��+�&���ؔ��>x�]�Q�r������e�aRJ�i��X��H�?����h ���@���c��ƛ���Y:A�0\�s� ���4Ǚ ���i�e�5�Fjj��T������B��C��W��o���v���?��W��;�5�ܼ�P�x�Y�����1��.�������󤬶a�$8>B�r�4����gHqIG#��6Ni�-Y�'f��6�%tB�T�}O����[��_�5X�q�BwU�49�e��) J��T�EX^W��g -��=�e�W�N�>[��JZ6�^t�g���̘/Q��Ι���A�26�ۭ]��M��_z�}tgݭ}H�6z�u(���I��2�G�{R���)�,���&�.�����Nz%�~E�V�o"��qS�U�4qɆY�&9I�L#�tTw����|Y��.�{�L� 0%R�Ba'�Qz )vJz#�������͚ba�u�[�{�~�8�L��b��荬:_�!w5/�����Tz�b@�?����$��F2_�s�V��kc�s} �B�C@��&����̬RזSW+�d*��UB#G�kc�4�o���b�Q�I���� �t�QHJ�ӛ�';��{�Y?��?���M�A��������0P�Jo���]����f�BF��I&��f;��-1����=�R�V\��JX���>���	FM���s�R�u���J	wnv%zbh�qrG53���`+����#ܼ�hQ~t��/b��L��O�3)XsWv7��1#{�ui�&�s70��z��> j3	�+��,;��h09O*��"����Lb��G["�z�*(H�(� ��V�"�*]���!�p�m�c`�n(O�bv��M���
�#�V-p]͒����	J�s��X��\|ϝ;�=�&�.R��ݠg��+�.��#4�<<�_��Ne�����%XLe�׋�[���OT!�#�S���z���ۑ֩z�;r���A7�t� �LA��&��E���s�|�{�b����?r��4��f�0Z�H'-�#E%nJ�I�[&U�5�A�I�@GiZQP
��%�^U�P�5FJ�ȉӦc��}��jRYa1^TJH��z5$��oi7�u��n$D��������dd��{�'�)X$R�"���+v��q�E
G��HqɽZ"u���p��Ssst��=;�FamzG����\�)a�*C��e`oF��"<�Q�=��(�f
�
��}Gu������K��9@�Uvi�찘
�����]�)i��H���֩N�k��AU3V�#U�� iST�w���q�^s���w6^^���Yx�ڄ�H�-Hk��*wK���$��	��O=�"�#O�vϟ6Z8�Ǳ�6��R?b�FX�yI���T
���Ec���C������������)Q��r)V5�]8U�iq���eN�˲�gT�iz	���g������J�3L��B�K�s��/�ݵ��wJwy��ȑ�X�	�!��K��#�.G~F"i̙]�e��Q#���f��48�� ����r]��BWI��Whc$'k��ľK�c3���V���0��cWz�r���z�IdP��XiM�?L~G?KhM�kAQБ�֫\C-L�kl""׵ˣc���Ьz�Lf{�~jh )�����Qb�aw������	�n{�_<P
z�u�E�d�᠂TQ����������l��CLL�5��-���5�������A���	� yz�"�4m��p35��F��I����1���/.����7Fz;���iw�g���0p�0��L2=!�ߞ�����d̴̪����b�L��6���ܘ�d!�(�V��&���hYJ0�Ω0�+�"�9b22�c�S���4��5��F�sJ֨��Z�w���jY�BHه6D��n!`���̓腨�Q����&xMML�*M��^��_�a@�J�+�]V�U���H����9w�wY��,"ۣ86?���|���m��/#5�j���T=���RGs�|:��'?�;�~ae�[�z��_�n��w�];�{NO �T���{�� �;���X �(a�Ȣ�	�
n��� ��1X
UW%I!��o}��c�Ri��""Ϙ��9@�;���61\�UX��ac�T"��;;:sy�g�j��Y�m[XS��)U�1a�Q���w`�N�*�[�r�]p*����ܽW�]ug18�(�O�� s�-�\��S�j��e���B�z�Ko���z����I/�D�X/�:�8��3�Y`�:x�=�}��h�(_�)酱Ѥ������x�m1�\����GN�2b1AzH,�)H��P�Ǣk�˘��X�V1�	}�y�Q����?����7�Ǳ�a��Y�2��U�- h#�b�
`h�0c�4%,�b�6h�Mj,�}��n���f$o`K,�z��¨2��[9s���i�
������I�͏0���g�4�܊t<��q��J=e�b)+�t]�f\�	�X����>�tl�@�Ru���ܚ����d�p�so&���\ �q�|�k�+����/�QC,�QYUhJII�#Ш4 B�U��*1"Gvix�6��\"]m�����j=�狹�xƗ�{�O��Qϋ��^����7K��{�I���
?�U�+��R���*I	q���K�puX�����L���c�}��Vؔ0�{���t�]�{?��o��ǃ��if��W�����>C㐓�9��Ǝ�<��n�ѕ �hm�P-�h\,�*ڄ����B��g.���_�U��(^��bh"���8��s�R�B��N�	ǱfO*�]*���{-M��������GR�܏�h�q i=�iW_�D���m�k�`�8���S��gT��m�`��p���o�]�$��Ltq�Z�4]�����?
,֚@[�ⴓ�Ü���| �53T���=�V��z�ɫ/κ& �wb�P�oJ�Y#JK]�l�=���* ��&�� i�.����$F���h^֠�%&-��H�Y�G9��>��Z��A��8�5��>��\q�4L�����50�w�>0k��#�-m9(8�"Y`�AX��(@u���Y��5����P��",�4ǝ!=�7�̾C,p�oc�M�Ż�$�Uǂ�"����ÿ��p6��
B��J�SA����<��ķ'S�k�0\s�K����1'���\2\���oQq5��1Rp��7 X-��[;�9ƣ��g06��9���K��Wݟ���'Ie�p�CJ�x�r��������8�����~�m���􀄿WH��@�3s��%����yV�q2�慕�*��0AZ5��կ�a���+\�c����V���Z�ЀV�؏/�G��c�W�����[�hQ�W^G�t)@��R�;+KT�1nr�'-�09��/��T��w��}�����}�yR�ϣAs������Y�q���&M�R�ٯ�/ �D/�S�iV���T�e���,oa3!�"�b=� c�����he`%�)�ʲ���{��>��O�WαI@���\�!��ʬ�_�{BBi$��Kz#1�RL9*�H��mJ�k��� Z:�*�Vu�[�cϱYI�m��*M<X)�����8eh]|������_	���*�m�$P��1�����f������-��S�4p2�T땆�!}���Oe`r�]��ѕ�X�O��g���߱���옟d�����T��yN�X]�U��}�Q-�?5~_�59��ah�4j��-S�`��Q'z�h�W-q� @��cQ����(z=�G���#x��	� ͻ?}�]�6���sv�k������^uo-lS/� ���7%49F+��RI�x�N��{l�O}q?�"��3A�5;L"U����bl5ᆖ�/��`�Z��� �1�Co%L�v�����U�G���K���c��D&3�X%Ҩ!L��C���ӎ�o�l3�l�>�L�v�JM���b�W�HL��舞$m�v���6�<N�k�FzH���:�!`��)�X�2�hV�ѯH�(P�fBo��}x���K�!���}=����"L����$������j�?�Ĕw��G�aUc,f�x̬�b4��9�$-�f���QEN��,l��}�w������0VcTb��Fnz����k��ev�89�HAD`���{�ʬ�N�H�e�Y�r,6G�<�vh�0�qH�9�xz�c�����W���C�$��2�^ܮ�C���P�R?ʋ0Y+|�,�_�L�_d�q뼷ʒ2{D|,f� e���#]3<��$�8��2����~�[�*�h�������r�%�?�Tn�%�u����`&`K��:���prin���p�5Oq~�\�����;������S���'>�TکM��3O�U%�¸�-�ƿ��G�~z�����- &����j��=�>(O*s�z�G݉3�Y��^�F�*�O�/)�� �5����U;�@���D�e��z����-�a-���P��Mv�X-|�h��}���{��S.Nܕ�z
W�&��Pbz[�D��?���d�����}�JM/=���>lvS-6��<\o����XAԋK�������YÙ��"5�_̻�s�?wv��ܖ_�cUBV`�k�џR>J�T��S��͕���,OL�_�=�E@A}���2^dQO�[0RH+��NN.ˀ���*c������X��m�_u{�����E]�E�2���#��& "EJ[Y5U�)��47�xʠǳ�|�%ur��،�DVs�6j*��E�]M�6w�}�����] �0)*���Z�aJ+���3�3N�  6εf]��^�,&FG,��#-|�6��ZR,���Uo?�ru�oGzem�Y:(c�����͇=���h�;w�u��k������h�z/�w>��޺͆�TX��_�D�� �����k|��N
h�x�x�Ae�ˍN��V��h���Tǝ���aЖv��U�׆	n���έ;����၁�_:0�{��X��|��]���
 ��T
�{��q�� ��3L�|oqx*�T��|rhCq*^���]��W5�|�����r��D���jukΨ�J$��aÊt�vkBhy�h����>!�)�.�ih������-�cT�~
��& @ �@�t��V�IT�%��U�KT.�Ӂ�˃_E?��Ο?�`��/�cG���|��L�M7w����]n @ 8���hW�E��%�]��� ��;�w�X��3��Am�W��O����ѹ��N�g����Ҝ�0�^Đ��PVN����3��~�Uk�?~��B�UR;j����������K�/ä����;����1��]��3����ZQ���g^���^\��g�fV���o�����aSHCɷ��7udFIا>w������|�j�)���x̌�&��,�/�"���N��u����?5�s�q�/���8G�\�x�O�"j4'�G�9k?��ҿ��:=ƵV;&�ǹ.QZ��ju�+7��D��B๡��e�W8�RS�� ��Z����3Tl)�%O5u�܀e�F��FK���#����P
j�c���H_5��J�	��o�����;w�0�L�lӺE~TUJ���HdO��M:����|O��#Z� J��"~iX�tu�k��_6X�K]��o�Y�*Á��P�_�kb*�Μ>���5��Bަ�Ňr4f��3�ro��*��uU)�(��@P�>+j D��R�b���ǬRذ|z�?Z	����@�U��8�����f�!�C��:.`�/[W�=YHcfoT(3H�%�e~�K���Ƃ���a`��x�`E��X�	��W�b; �&���xh |b�U�i���X�̓+�����2�K����*.Xlq�@�?)���L���^]�y�`:'��(�W��
�7ZU��c/*״�?��g��	��`�Ӹ���:����޿r۽wy�]Y߅œ�+L��O��l�☝
����ii]x��d����8n�+�v{�Y�<":�kT&{����LVr��.�ʖj�I��,!.�n�Һ�i�Zإz<��GW����;�qd��G&����K�7<�nI��"��}�L\�#A�8_ A'�����і��v��]+��7.��P�K��(�@���$*wn V�c�\���1N#�*`��v�-D=T���B�S`�L��g�j�:	�Py���Fa��ـՙG73��IU;�<7�샾Tݔ��_�����M��lX��B����ֺ%�%6M3M"�^��S��v��O�ә}��>�b#����h��~��ث̚m��D���>���Mh�����K����X�Ľ�m/��Q�k ����c�w�RQ���y��}ī�BQaҤz�槯P�S��g�}��FH��QY����#[ɹg܋� ���G�0N<J
��Pv����y����Pe&]f0�x�a�G�t���=��e��,ڋ�ϯ���P��f���@]cbo����	ۖ����h�� �ѻ�J��U��ھHl���+���%R��#��E۵ʢ�桫\w�?��-R�?
(�N���B��$��b_����L�FI�A�uo��G�����!��
���Icjq���w��W� -+��7ga~�� �>�KZHk|�޺i��} 5]�D	�� 0`e�)+�Z�n�--�%�S�N��>���V�z�)�;J
1�xo�.5��т��H ��z9�k���;����k|°�© �N<Ú`��ϽVg�/Di��y'YX�T&�h��SB�f4h�{�1���>r͍��	���Ir�yQ?/�v �hA�=)z��k�A�:�����*�6�F%�����x��e�*��&� �ʿa�ԫ���gb>UI&�'ѹ170|{�eVxabm�ǋM��X�g����T�5`�X���Ҍ^�m������2!���5K�@n\��I, �HJ����DD�����H5�Qbbb���-*�ȵ���%�������Q0�--#^+p<Gu� ��H�d�`�)}� ��9y����.1t߼���a�H�Ȳg
 �X��w�0{�����9wi��>����k\GL@�W�y(�
��ՔN3M���>��8��A{���PQCV����IC�����%ŃV:r���H��b<9�&#▘��=#K�o.�����<��щuki��т��wT��MԚ��טt� �E�$�H�%��B�L�*��$$�3460k[%w ��x�=�3�Swx:���9^8�]�x��	E�xg��`�;@ڣ��i��Xu��B�I�{�w���ۤ,�n�L"C|mx�$i�d߈[���945'�6�g�TP��D�Bo-��D~R�a����|��Z��0H1<t4��5�o��o�i��;��M��s8�ʹi� �w��}�+�L�a�]���"Y����O�>��_�T\��c�C���[_"��Ix�.�s�H��{�)e��<K#���a���L����)�*��vk������(ᾆ�䅗�2p��`ez�S)u�y7�T���������Q?�6;vU����+��H��Sa���o_t7�� $Ҥ�ڤ�� ]D��?x�=��\����["q��c}���,ܦ�N�k�2���&6_H�SF��wE�<�1���G\	J�wamVǯ�G9�� �1��2X��斻F�7H�i�:r<��Fh��{�����9#���u�Uz�����D�A�J	��JF�k8{�i1na�	4>8L�L�*�a{
�L�~--d��D�E�N������G�wܷ_��5�=��)w3K�5��(c����i��D`K�ɱ5Ͷ�h�8��?{��di�fgb۵�Z��#ufUeVuu��j	t0��9F���xC����n��K����ԙ����p�Z��~ܝ��~��\��UdTyF���s>����^�z�j�o�Wj��OÁ%�����h�b�2N����-��+4Ip'�&�p:D!�B��"�� 
0����b��*�P��{5��ż���x�� �.���`Z�i��N0n^���Ϥ��bo]�wKh���5 �c֘�7���2T2+���-��nqo/�)�j�s�PM����0{�6aU��9?V����˺ع�������.�a�(�	���F6�G,��&[���.H� S����� ��k��p�{mi�f�">�13����Ay��u���V}޿B�yK�p�L��q��B�
ߛ�s�8lq��s�8����j
gq�pY(��/+���!����X6>�O� =��7|}������t�(�)X@�?k9��&��Kq\e����҈�EB�������+�;�h�-�W֍��%SX�`2�)v�3������d<-��WV�_ށ)О�E�u� ��z~s�����_ܛZik���L�xw���J��LPR��'x\e�u�Jwe�Z�C�� )�-Ҿ��Q�h� �Y4˘����'���>v�̢i�����ؓGi}�������`?�  �)Z-@�����bo����xx�h
�t�-l��y P%��3Ц�;0 U ��<���ȱR3�IIG��y|e�jbQ�⼖�Y\rL�Ի���K���gY�Ì�X�z�9��K���|o<��K�j����7��	�ɂ��-�4d[���'�&�K��1ϱ���s�%�~�����5t�tx�T�Xm錅��矇����>I�wn�b;w�F�aa6z��S��E[y%�����W�bA0��`
��$�m���ｗ>�3�2����49@�-�����`��D�|)����K��OOGB}�9k
�)�\�������x����_�[���c���ߥM���4�;4�<s��FJm,[0Ni��x4����"b�FDɟ�'TU���MZ�M-e�]�ke�C/>;�*���[hkR,�a�O(U��Oҽx��d�Xe!`\���b��@����~�����'��/���ͦ��}�eZ���"��>�c���1v��y�De��]@P l`�cS���!�i��%�S��uc/`)���
@WuS-Z���˿�~*.�#����<��7h�ܚ�lV �%h�c1��QI�;���	��J�:�%-l,°��DV�`�T?'��8�,k��.��׽:���0���^Q�[��.-X���We������-5��m ����u�F���b�}�4�U� K��68�2�1W\g�R�b���ˌ?��t��������9�!�.�d|W$EǙ	��e�/��a�+`�Cvu���=	F6{{����ej�X�#Ėkm��`:	���PGݤw�02-[Y��܏�F=%�*�q���ܰ��`�|E��k<�2g@�]�*0��s̪��lj���l9����e�T���`̧U��RV������p]f��"���ZU:�_�Z�1�[�����(3x�+��8��S����@�$��i���x����tv�r=��{�޻�V���s�	�Ջ�L=�|G��N2�_��"���<r3���@�w�ѹ�_w1�b7u���w����D����Y����灴CjM���T_m�ZOW�ܩ��U|Yj�ۛ{{ۚ[�+k�ȶ
�m�ur���4�J��B{�]�g��"6Y��4��1�;rx$��g�>���~Q[��������vs--��"Bu�U�FB�C�����_j��_$~�	B�6��vLup� �{�tUHxD	� �ĩ��T���Ȗ8)_5�f`��� 82�!M�Uܝ4��Z��4|�'ve?���hU�� ��ζt�ԇ��*��,�ݰ:��8I��{�O�����>�ҝv�o�%�k�4yE�vm;w/��ǅ�����s/��s/��<�Ϲ�FgB	�3Jo�~��t�pY��Z:�8��\k[��I�o���A�k����Ӈ�L�O�
�w�E��E��]e�������x��:u�����ϥ��u�}0�t��N��B�%���Ֆ�+�%Y� (|~�G?�E�����C��Pq�4~,V�-%���i�E���/}�`c*F�5�6g����ҟ��v��y��z��I"]��H�A<��_F%`)H�=�E��ԫ�����0bM��eܚ�z?�����8c�ʱ���t&�:-�BMs>/��Rjc�}�.f���uʃc�G^W-�Ǒ�Φz�'#Hp=�6I������I�s�Xmԃ�<��:�a!�f=����;�?��{%���[ߠ<֔�Z� 3��*ƥ�L�}ّ�����Xī������(��fn����2 ���k��7֔Eg�M��� ৱM���+��[�."����ܓs6N���T��̬���\9ǥ�P��`�dÁ����X�~AfD��b�;2��Xz��2��)(0��­���-M��(�9	N��Hˀ�m����>�3�0F:GW	��%�]��:�zA��(����!��=�E�^��P�q+@�AP,�V胊zE�,!k��X�-���Ua�Q�3�X����J��U�����Q ����F�d��\?=���{z-��������,�.���)1�7��N�:�'��d����9;�eϾǟ�W�`Jwk�xr1��^�>��c3i���T�22J�\?Cn7�����زR�!�?�a7@E4�c���^��y$�ɘ=�����vF E��:����W�E1a��E��<S6J�Q��ML5��D���v���b�c���*~*���ä�v6!n��K�w�jjXH5c�gUt=���Ҙ]Pt�t��S��oz8���Uf/�� �]�?1�c��Iڠ�:vq1��PkΎ�%0L��5�����Q~�f�U�:ǲHK��5%��c�6U�FR�a��b���u�0�5?�S�s���ZMq�2K�q�RΔm��Q���;�@�a/�{t�}���i0u�؈{����2&�\F~���uu,�V%,�=�;�V2y�zZ���bR��7��܄\sF�N� �>��AK,N[�����u������/O6����#��:45u�p���aS��3����zګ�)�-��}�V�%4S���{��G��"@�d�� @ G��Д&_P������g�[;���w��`�Ǆr�2ںF��3���\��vQ���h��1�q4����פz�L9�b���Ѥ��@�dmq�p%[��/l��X*0\�$v�7��b�E��<�Y�N�y�`���.�RJ�᳚h���8���=v�sDl�z��4:5�6�,�ۈ�?����0��^A��X��0Z�&�j;,�k,|���,�.2�Ս��jYΑ%*�|��E�pU����\���?䞣E���,� e�.�QۂU�S�]6e�=��胢�2�`�� ����Sf�4Ю_�5v��f3��K6�_]�	m�&���m�`��`��W�1vw�ai�R_����#�Q��u}�M����"�@n�����o��U����e� Y'���ܕ����x�Bg�Y�p]��55f��9s\8��9���1nG�9ʋ�i��$�_�e/,�[��z����TEƢ�m��b�p���}��d7V�m��x�lS���ҙ,�1Xn�b��e��/��㣣�L�+c��jx��K�'��D���6�I\X��UȈ��S�]b�/����ϖ��Z�料� h�����/����ׄ%%����߁OI0Cٚ�1L=>�h�@��pz5]�h=M� �V�m��S�Y�F1�8�w���pۜ�&Z DM ���s-���;�/<��;�p:�/@s0)d�A��~���	*3�*eb���O�;:�c�Z�����c��W%����N���\�b�j�o�s;�uʹ|[��	L��g��s�C���q�C�K�WQ���N�w�W��\a(�`g*iw������o�N�_�, U/�NZ��`[h��`�n��QC9��k1��27�,R ;1J�`��F�ȵa��g[X+X�a"�G�:c�JG�
��	�0�d��
]�;�u�m	�fCP��Z!���-�#��G�\����N<z*��#��/�O�Gly�����ȁ�B|���m�	�g8�nq��玧��#��WR	���}A-�PL��7(�܆�Y��������f��Q ��s˥yv��h���q��UEG�h8�Ǖ��WY�?f��1��RU-><��wp�GHK�$�g�{�pSuz�<��d�maS����-��?�mz�_����b1�[ci�C�����9���0b�^ �k�N<�M�A����D��÷���� u=�v�R�-x�L9(��ߌ�{���K���6}JgU���A) y��>��E�7ז������e���	e�1����oCԬ�c��}����븯g_{5س��S���^�H��T
��=�s�w��>�h��э;i�A����b ݒ�.�͞����%G�b��L]\�76�� h/��Z:{�t��s���?#>�����)kE�+�Bp,b���J ��s��O7c��-� ����6	.��h���=��\[I�1Bm�:������H�t`_�{�7�8�n�Os���@r�+��ۤ�E5F�6<�מ!����Mfj�����F�M�y�EۍC�.�>�t�)vv�<丈��a�g�/ S���P�箏�Ē32,��w8�KVjNx[���ir"�ݎ) �.�E74���%	�2��,)�V�Tn�s���{ع�s[T�M���R4aS������!Z���li9��?�<-	@+��.n\dB�F��EȲ=�]�0c��۲Gv�Hq�꟨�1wm�i6s��1��y����q�������,<J�Uv�r��I�Ǹ�`�H��e�y|���y/�x�@>E�Y��oh�*8N֝�3�R$/�Q{�E�i�V0E��~�+�_��AP�iZf;��[V��θ3�Ia��iz�n+�[��`4����u���ke����#Em�����&� k<�;z`�:>�Fi�'e����E'޿���Z��'w5�!�0ꋽ-��\:ک4��F8��li�W�}~9�MsQ�Ȩ�
��v���1�v���!����i���Ew�R�Tzq�p|ʹ�7� .��V�p�䩨㯱�)��Wa')�0X��)Tt�7�f�������ϋ�-NG�4��*�(���E��V�� m��X�>�z�R���B�M9L�Y\NEWC��O/�;�G�}
�hA񓎞;��H��kj]U��+]|�>���i:�`@��x׬�,���/�+�}'-�Ҵ��>B
{+�U�Q-`�K5Z��J�wx�,�RϟEp-wiՈ�W׈���r} ��$�WpӲ=H��>f;@�j~�Ż�(��˔�kY��>Hs����R��ܠ�Ŷ�=@ӡS�RQ!�G(���D��Η:}h8�.�F1K��H��{ ����]Bi�&o��-G�mLX-��(���ɵ��m��\��V���K���m
1�: �� �Va:�Y������NRj��W�M�L6�>�q)Cg4��mI�o��&��M����t�a�@��]'��	Z�G^�mн�k`��s%�v���}��a1���i�::�f�[V�ٳ�*@�ϕ��N�R���>�:O�pmU�h��ҧ�A����U����n���N=��=Q��B�A3Z��Y�d%��m��a���,��SvE��EY�����5�}��W)�m#���r��זn�g��^!����u4���k��7�pF��.��F�q,b���~7�\aۻ�f�����@dl�Yc��ß��]�j�O�<;!w�A�瞕����;��������=b���R�^��н��F��,u�~a�-���dL�,�A��sJ��9fb���(�3�c�.E�e,��9�f��rƸ�Zv�����|�0�q��Z9��7��= �,�Z __
 ����UC��=�^#uB�`;�M���J��͎��[+l`��SZ��<�v��*;�
�-YE'���#�Ɖl2>������}̕������X���=�gʴ�� �[4+�~:aGS� ���+�_E]��__�x.@;�v���<�XȞȌ�1���t�T��]&�[.��p���f�D���:�r��7��B"��IC���u{d����R��GE�c>�*�4�L w9]��o��ŵ�;,�}@������?�1���Pi��;��	��)E$�)b�;a_�e��ZGȼ��U�4�����H����\�Σ��ɵ�]�;H�t�� �c~']-��W1J���@̡C���#�;�V�Ҵ!�\��IDʿ�����H�_����Eù������BVj�]g���i��(���`Z:Ky�����"�ή�EG(�����(���	r6�>G+wå�`} 켟�M�?�<����Ԫ��Ji����3��q��
�s���	xj�L��x�����6{e�2�?������ ��)��Q�_W쎾��O�����"ګ�S3��U�?���#ڣ��"�{L�� �}��#�oySy�{N]�\�gRs#~7L�� W���~����ǈb����'��H�x�����u��qO���>L�J�C5a�x�qL���+\�&���*!qˁ�4CI���5����O��J����G��s������s��X�d����h�w�>��v�q�GS��;�O�{���!�w1�m�`�� ��-��h�Pq��N�xn�nJo����	 �_���񗦯��r��m�r�3F��e�6�L����,��i���X�ݍSzcl���O>Imt�G9���7��"����]f��Jߨ�.�A�4%Ⱦ�NC�X  ��W������+���`�Y�5�� b��+hi�&(J6�%�8��.
�u\d�E@f� �R�Y^�eƂ�Pj�,�����B�N�d3�\X%,�?S��x�P��ka@�� J�N
�y���T�$�c)�Y� �j':�,}9���Xr�ٍ�(�g ��O�{fi=·c��`����F�ܶ��7՘:'�i�~����sM�)Y�U)|�@(������JMh;u�V����}�;dx���r�o�4��Ŗ�R�&��1�B��1{xĵ�Q��������7H�W�\���9��K������L�$H7�����^��� `%�	������u��9��,���p�:�֝��1&��m�ð�3��|���}�xȲI(�䰆��l�y�?/�������v:K�S����Z�1Q�K�G.�c�l]�M�V�S�n���i�z��ЅTᨙ���yΎ�3ѥP�Mߓrg7^���B����q��P�����)��'�-�ˠDr1v�P�Ao�쌺P��~���1�6�V��_���E����ND�[;���g�{�|̮��Zv�y�U��
.�+��z���%x��a�����6�5�F'�ɇ�i�F]�EsS� X�����,����N�E��1�kϥ*�v�u��n}~%=�Bxf�Pڇ��Aq�����������HNՙo���c̈�g�E��� J�'���?�(�Cm�K�a�KH�\ٌ(���sv�=_�M/�=�r4���Ĳ�/�
�t~��� 6{�cp����s��
�e U0���re�7[;F0�#~$�%�nӴ�07w�_K����Y���q�wє�]�)~�]ZP_NX��8��s1���2�7�[&���ie�1�������=�\؅�g�./Kw�o1���z:30M�l:O���-��{v�y�;a#�-��9ɎX�]D�?ׇ��f6�]��G?'��G?J�a�:`ƪ�sB�{%�DLT�`�\3#��Qt��lDo�Θ�7Ic�J���"����1���w|�5J��M���xV���z����;�?���R��v�=(m�A��PR��-s�Ŀ��a��u�+�$�0:l��	t��(���.0�H�Z���zj%3V[�#�>�U�� YQ�y`�9�Ke�N�9��3��j��Sv	.�yX�5;�b���M �`a�X�#�D&�.+���F���w"���pj�輚��I�R��q]�|d��r�E%�J	Q��</��̕�eх�1׈̈́$�?g'����$h�)�IhN��_FiJ-�`y��w�[��U=�;ʈv�1�ǹ�Ѭ뇠���1�L@�誋cd}Pd����h�/j��>�9�@&kR\�g��/<��\� V1j�����P¬���bRP? ���Lr�`�u��ӥU7Zw7@�x�Bs��5=4ni&H,e�Nl����!U�����ﺠ�B]��p���')�t{P�b`M}�ϛ��y����sF (Z��|昸(����г<��� ;:�?v?N]NV�ѕ�*���b�?L�I���!�����@�և#Dn���#R��dIFm_�aS8��)�`�A��7w�<1{E)�rU7��}#j�3��8Ory]�F��ޣ�
`:��f�i��ޞ����Q�jEP{O��S�i 9<�R�J��<ǱF�����t�4Qj##����oܢU�n,:�z����|<s2c�ہ��$��C��HE���8��>� `W�:9_i�}~n�ɫg��#G��g�����;�˖�#u��w���DO���i@ ,���Te�eX%E�-8.w�M������I[m�mT���_���� i�4����u9<q,��LD��1��WWKH�4q�\�.@Ƌ/���p1M�Z���bb�i�I�?��)$�e����9�.�Ri�_X�3
���r��NgTb�ğeܧF�YYG# �!�}��Г�(�Q�z�����0pK��߈����^M��j���s�SJG�:��[:~�!N^�� P\�'�HU���r6:�ۅg�
�E����~��������(�5�����Z��A�0/+��xN��V��T-�"�xBx6* �:h�)Vj^�Z��Z��폋p�{c'�*��L�û7�m��Ry�Q}�鏿~�{��.O�*�62ƲEn;�@ +���!�����PR/�� �gR�rEϊ�m>ȗ�`*�u��o����n>���#�=��^�����P�Fȹ)+%�D��Îs�:�v�&���A�e�s!M8�[vE7�ˀբ���
 ���|,��R��������_̥��τ1�lX�c2ې};��.:�3nm��2"s`0O�Vp$�c�D�s��+�5SSS�ZZ&���y���J�ez,3�O��3�y���OV�3S�ǁ�l�W�X(��}z��g��3���U�!wlq��N7q0N<� Q�?���:�@gF��4��>(E<װ�=�����#M@�Đ�ճ�0�Wg���k.�;���;�x�m�� o_/!if�1��#�1��:Z(k{�W��t��<&������A�d����婛�"�X����4=���� K9L��Rt̵t�.V��	�=��2��A��%L.���g�ե����p���T��_cq�Ӥ��?�g2��-0!�sw�h�}�]� �I�ҁ?�낪볠��`4&������躚o']�l����8,�~�)øp�pZd�9r��'� ���Y ���ُ�y{}��'��Ŵ	��E�����]�a����rJ;�X������Yd7�ѹ+q�䞮>ڝ�S+��J�<;��?g������#4,i��s��>��~����"��-��A��ꂕ��ld2c�$��q>5�L��	6gX�=����ӝ�wҝ˟����X����Sޫ
�:�6H	�(؊Rʉ���-��ɛ�c7�j ���Ͱ�~�q��l�ѣi�jM�z�}�x�R�<,�2�a��.?s��Y�׸������C��̹��%��>���m�I����ܸt	Q�p����1P�1Z����H\#������v�Uؕ�N������!V�9�;	ד�k*H���5sA�M�8Zk�)��W�{��M�^��� �6� ��c:x��|k`���{= tlm,ݺq�ԓ��f�-�i�g���E9�-�U�}��>�2!���{m��>$�M�G5��}ƶ:�m��`g�`�v i�0_V�&��o�v�n����4�ӔnO!�e\������0~�و�����ev��ܣj�Q�\�N��m��@� �v�WXt�𚱔��t9���-�e�r\���\�A秃����X����M�"3�-�l%�+�͟��"�g3��.� ��> #J��ѱ9+�G��J�X��\��v�ɴ[�۬;,Jj1_��a�㦨1�v�A�n3:�3~�. �'�B8��F��6|�,Sikg, h��p�~dq��n�~�=�]�KR���Ni	gI�,2�t�V�����9��2=;��a�a������D�s����=����M�!��5���~�=g�6ʅ��4�� ����� ո�%%���?����c�
���#��lF{�s��> � E���;��>$p�<x�j`ad�L�Y�Cv+~;�I�S*e�`��Pg]�gw=��ݸ����q[��ɺL7�)��J�`��J��ľ	x@4ډ�N��/f�1;��=�Q���ŗc��
tI&N#����<z�F<�-����u�I���w�.���d-�Z����DYT�.�I�aLD�#IJ�%%u1�o�c�}�J�r�}�QeRX�kf���b~_��$^��d�{�X�'Hu~���}�_����}�d�E   IDAT�2ܽ�i҉�ֈ�t��u���J}[��	f�i�����M��wX��)�=$@Չ�$�&?��ۡ�j����zKVM�[(����sV���7�^2��F��p�������M������V��0,S��;��aJ<�5��i�u�
�T�y����R:zH��2��f�;�ek�]��(��Ꚗ�y���s��8���0~���n��� ats:�=]���M+x"��?�>��@���ݽ}l8�vo_�J�:��R��[��L�ߑQ'���3���V�V��m�������/-#b�����2=��{����-.������� �nJVy�e݌�l*�����6��	4_O�3�s�k~b,JO[��~ޣ�hlJ�D0�� P�1���p�O���袚{��~�W�����hX��g�m�v {,��j�����g�硅.�G�U��u�VG�,�z�wP�������D_vo�
ʈ#�� ��kΒ�vg��#��F���E��l�:;�W,�e p�(�y��{=�fi	h�i�\S��3KC����G��vM��r�JJ~�.b[R����E߮#�qBse���l0�"�C	�$�s\^�E�FѰ_$ D{�-{:G{��h��G#��d��O$��e��!�i5�� 	6��1�C�\p#�r�7(|�M#� ʷU��x^|��G6�Z�-��a��	����W~���~��R�{������c7�m@��'��m;�u��Ȥ������$k˜�,�����6Ƕ�G�6�����������3�e|�9iQ�K|�/a�|�&�V�Mv��~T��t�y>�G����h�s��]m=� h�SV��e�j�� #�,�UL��<�U��nS3��E��2G��H
ReK�3WC�����Ig�@w-�m�D��Y����N�	JMcD@��Q�hl|}eE�S�3�e'� v�w��MA��;�e��3����P%��s�[7ш�&��.(��}��Ҧ�?����B���/�n��?��Fq���p��W���5R^z�H)m3:~�p�^^��#<n���fT�
,MΧu�PW�ӯ�4e�I��s���KO�ߊA��%^���\�f�] �b��w��\�|r�J{��I���z���:آC��/Y�y��}װ�`��&�����tsl���w @��!��ۥ�(���:`Ǝ_xg�| *����;t6�~���?L��Ͳ#�}�-�V��)����9���$#��N����b29���c8� �A���ݿ�f����>���9�����8�jA/�NO�Vخ>�����}�r��:y@�}��l��g逡٢T8v���������J_ G�s���s����v�vI�fL�ǐQ����<"�qƞ�;�y�{��׏�/�_� ���#tX�=��AY�YH�Q�-.�ΰ�W�S��D�s�< �T�a|�!&�y��u���a���Y��r�q��/b��c���)�]Z%�������c�s�=?��u�"鯤f����#J[00��!�����TP:U�����'���l2�)ˮb��HG]Y�W�1;���^Ճ����U-EuP�����HKu)�6mm����t��uRp-�������_{	�r@���1E�G��Z�Z |-V{�?�m<�(���) ȭl�q�a�xD��<7݀�F�;�k�[�.Ԕ���.بq`�QKlx� �͞J�8g(A�lw��}���-����)$fv"�n��v !Y���`~�&�����K2�Y2��H�!�d�uB��	+�LE�!�Vc'h�ˌ\@I6� xMA��U�#]S�=���*��U|�%;�F;t�k�8���y�I���m3_�U�昻�d����>��S@�6�ͭ҂���N��dhKC���a�Q-v3Ѷm��$Y@6b�{�X���3��Ke�� ��+PVV�A�&����Ta�.�lǃf`�|p(,�Aܕ�l�0��������P�@�!_(�˺*��*�"��ePo���2Bϲ��� {R��Բ��f��N�ȱbg�	���%8��w�fǻ
����|���&��N�uz�b�*Lf�wB��yf�umg��uZ�W�6�q!c�k��K���%�w��Tl������ٮ1!@�*&����8�J3Oa��6HG߽zat!=���i�Ko��F�b���
k�ٗ_ �j$��|���+8��t���4�����:�%���s�֘,�j�uc�G�>��鷾�&
�Ig��?�_mCU�v�3Ŀ�0<�I��&F�Β[�P�i�/C�c����VBWF;���
ۀ�1�m�X�i���G��N���N�I�\�Z4<^�}�X�},̃a�g��������i�{�8-?��P���G�}�~�W��1�M�Ð�<5h
�v~�n�Nr���h4�3JGޣ5�0�)=bAo�]聉z����Gz�c�kc�W9cB}���v��:�h�'���.P��0Ja���0�!�eǧ)�^����͹4�}�a����3g��`�,�G��"�sr-�1���/��^ۻ��u���<�a3_x1M"�?��g|���d�O����<x�>��;����}/]|��c+5�no9�����3�{oS;e϶x���f=�s'���i\�e�b���g��bz�ko��!��;����b�\=%�e��&,�I���z��F²^�Vb[��{Z����Xl	L��!�����-��5޳P��{mp����C�
Q��������bg����'Y%J���eS@��3@�̖l�Qy�MK	�^����.�	�>���k٠{=ƌ��z�Sç9��4�4F�G�2�m)�2"E���iժ~(Z��9�"��ι�v�%NΙژ�F[�յ�N0�j.굜Sޒl���M���^Gj��8A���Dxw�Q�p�a�h���R!�2��lzh���|l�Ǎ���L;�;k�{�j	+i�� #JY����ʧ�7��v��B+ſs����Ϻ�Z�j�u������%�c�V�0���x	�v��2.<�
X�^�FuKk�Je�S�?kԧ)\���6	���,��Ѻ���:��;��_��	�����;2��A��+p7 �| �S�c�_��ï�M��y�ptU7DwQT��h��>N�ֆ��������.0�7񼰋c����=��-T� ����8@G1������ח��5z�4���N� ��fX�=X�[�����+��yF�������i;RK[�fi;�F�-,6jy<�ؓy|v�S����@��;F��Y�C�
0�!7ɅV['�������٩��UF����ı�g��j���l��xzO�? �Щ�r��	�.@ć���Nz�+���}��`(�h���Eۡ. ���1&����,\Ӕdn�Y^Wn�L�������=��?.�𴠝�X� /v���b��\�GNY�ݥ��?�wd�,p7���k�_�z�Y�P/	�G�n�F��>I�Z�*��-�Y8G	��_�1M)����,�-��ӯ\��!�l!X�^��<���9m>GjA��ͫ��fP���͏���A=���Hy"Kz�ǽn�x�*���IU��+��p���l�{U�v
���zec�>N������j��Sv��h��g�e|a�47ld<.�.��s=J����Q�YCv6�(�4�1\��k������.�,��c�t��X��@3�u�kX��NE�I��$˵�Cˌ�-�@e\kw�K�\S5$g��L�#��7�
PDg5e��Z<�7d4'��0��n�+�V�&꠽��F���V o�K`�rF%�V���{��7Q����)g�ͯ�MÂh=�k㔴�5˹�Bp`[��a���\F��ƣ��<��:L��ř4Oi9O'e�5���"��vu��V�u�Q��V�"�s81��23��a�4��am�t2ח�|��Y�˲�o�^=K���.,�-7��t�� ��i.w)�e�o�i���W ���D�h&�6ę1��C�:\���+Q<nW]��2���e_u���k>Jk��~f5P�Y �e���}���i��ˍy���Jn�K�-�|H�A�؜�=v�{F2�g&��K�W�NA c��K��ca��|�W�� A��=�>G�w��q�	:b�?Mə�T6X�#���&\��������XwQ�#��d��&I#�`�����#��Saq�u�����!�Y �4t�N���eګ$CC�_2A3P���2���p�! T�}�f:�Qd�o��ksDŏ�j�*�^��t�����~�4�a��;�f���e9Jqo�+bb�ϰ�� x�py�����S����(=�%�S�]ϕ=J#W���|��A���$y+xmDW4L�T%;�~ N��cJ#��Xͳ�^a�_�E�sb*]��V:�����4Q������3�(�m�eI��ϧ�x�y���~��%���N�=�]#e�z�y�!�2_��?I#��f���\�֑�t��,ۛ���ӊ3M��]Q�!�9�t��PR��w��ke1|�d������6 ��2�^\�����/a���
0�>�w���i��FSC���Zg�ު/O/��?O���[i�Z �]xtq5�Z�q�~��r��V�Ey���UF�m�k�dj&2���ϱK�Ko'@�L�,�>��}}�K��&Be&x�K�>���K>��cܟ��|�3��Ʈ\��U����շ��n dv|�qU�����çi��,Z�U�)��'p�>q4�s(��z:/#�������506�p}
&m�q����4���q����H5��,���ճ����e&���K�����%���ϣ��"č��<�p�le5��M��}�>�]@�R0[�&��#S��_�t
F�es=+��w������Zf�)��D[����mu�M���H�/!^g;��?�Y�T�YNr��y~Q���U���T�ݤ��SR�m��?��ք�뿦�_]��w���~��`�����s���X<�R��wv`�u�^ ,V3���N8D�nGj}�z� ��Y�,���U�_qTzY�r�O^�"�A�(�v�u�E����S ��|���]dt��h�q�/5A��+�Y�$Y�r�D��=.]���动���<����v�@t��S�6���2��
V9��z)'��(p����5���{�S`m5��rFV
�E�(��Z���a��F�,56���c �p���w�ă8'X�y�̯b7��ʠ�vl�z��B����	I��҇܇_�.�j��E��ur۶E�!�տ;�,�����d���ypC��NG�60-�
�c������>	��I�]R��F"��g�.�x �3�?�ʴ!�N4F�I�O5�h�w0��?��OYT�����I/�2M��3G6H���S������h�㩧p�� ��t@1K7��2gϞC;ѐJ�ʘw��2į�=-��c�ZL0RU,"ˀ����|�hE�/��l4q�U,J:��^<��1���>-񞫀�vr���F���_��i�X30�Ɵ�%,�2:��DR|3:��ޣ����V�H��2e�P_7����?D���0��q� T'�-&ԡ��	Q�g�Î���R��2��!B�q�ؽF��`^n��	��'�]h�4�5px(ʬmx�=׹��cC�&k��!�hP��H�v=����V��km�\A��Yg#��ة�6�*z�;��b�`IN���nV����Տ�P"�=��(������E��o�+&\XB���U�I^ ����7�� ]�s42l�F5H��b��$%ū���<�`M�A{��@�Ϊ����MC�|��;�+9�����t��,sA��s�����:�p�Y�uQ[�u��F�,v��Z6��[����o��Z��_�f�:e���z�$��ݝ� B�8tw��)���b��u�!���Չ�h������|d�,��o�1@�la��:�%��7X�g`�Q?#��,�~�Ё�Q��3��U9݄��|��/��"�.D��lB}]�(�x=�,_t"��3�5|�ٌ�y��$T���m��=u9<ky����k����a,�������ۧcͺ�=Vn�B[㦎ۍ�rq�d|�ӥ7�f*��|�k��)YZ��ɚ��GMbnYu٥��.Q3���+��!u`�?��D��m�~�x���sl2^���\�}��gZ,�"tKm�7�1	�4�<C̮����Z�C�k�p�V
�,#z���]W���l�����oԐ��E�N��O���g@����%�	�Y�Ut@&�c�:�V��������Oz.@����L �Q�K���j[�	�g~>���x�0A����^m���)w�!��	��a3H�2�t��[j4���Vm�;��.:�N�u��ڽ�7a�2�%�4/w�!��t��2R��	J>���Z�sk�!莣<��p�S������Svv�l�XO9Zz���ܽs7��������r�z:S�����i�-�Y�#�!)�D��0����;��[Y�+����$`xfY���0�	a�k��CtM�D�}��n�A����x
�Cr�����u2�jS��&��5�e��gGo^����:�^Kd�����"��`kj�����r�}~�4r������3t�T�ҩ�GY�
87Ƶ��L?!� ������]&��/�OU���<̀�m�>B�ً��m���HfoM# �
�;:��X����ƍ+�(ᯃ�Ì��Y,�9�ؘ���&�	�!�X���qc�h�~�x� �V��3�)]K{�� ?���sR8-�۟$���M;�����_(�7��w����Y��+D� 	B�"F�7�~�o~��?�,R�-��p�('��w�ɻFF�f�:�A'LU������)�1"�͘�I��"�Z�o��������}͸zߥ�v��Oh'oN�� �������{0\q�^ܹ!�0���Tb��"L��f[��h���sye�9D�M�7y�����ƈ\y�g��	:����I���JK�G	j�5T4��o�Ĝ0�9�}�&�Ȏe|����� G�҈�m���U[ᑴ)��1��a�����ۆ(�"JOf�+��_.�<O��5j�ؕl���x�k5�ONK�:�������D�F�g��r�f��������V�̂�j�Q�k��� 'q�"��}���z�Xj_,��8�a�@�l��1_���b@��df�?��2�14-XV�����Aς��D'.��ne�5#tC��w~����D�,ۮ�fҼFI�w�X(i���55Avr��2�]�ʿyN��'�Ƕ�����RۮB �T�@dW|vh�8;�=�T��5З�NК�yո�̀q0[�ـ�������/3^KRgCM�mes�=ycy��k��8s�!�;��ww1�ei�z����|a� A����K�H]���ߑ�̨��jp� 5���6�ѭ�~�����B6���t�X���y�4Ϋ�vr�x�������iA��v:�t��Cu�P�Wl�����2��]?�
�mP��~��Xv�PX��>�2��{�����s�ѻLd9t��<�ۈ�/�`��@�c��@��� ��8 F����w��-,
�,▶��j��B9��O;"k�\�ж�ɜB�5v��T�Cr/��K��(aT3I����o�\={@�>�*�����(_���&��x�.���	���]';���*�
�^�Jz��~j��h��N n�g�/�3^�����[��?  U���� ��3��7�:I]?���	&���L�k7�b8\L~��?NO=�:��jz<��9v�w	�4v�y�;�=O����O���۷R����X:1r<�p�B��/�I�^��0$��W'��ˢ�qT1�.��1�ə���o���V���;�=I�-W+�p�����&6�E���wS��Ȳ����f�u��X���5-V.�z�p�Y*a���n���G�� ��V�0���t@��uSo�f���@Y�Vych`�KX����>��	�U� �"�i腳�����7�8��9��f�7�F��';N���#kN VI�����ͫ�R3b�^�S�;�� '��R���Ǖ\��ߓ��x0G��<1�Z�M/�{t�ݹ~=�8F\b�2��e��rY[�Ҝ!����DB���M�᷎��jʚ�A�N<ET�۲l]e����SN�Z�q/��#=��Ӆ��Ql�˜�b)K���< ��yl9�1�@ld`� $O�F5m�����㔖5�c�s�����ۆ�~tn����.ږ�X���ÐR"R쨂iܴ��q�HA
�\`Tm���5^O3�F��^�3��6�Y�<�[P[f�k�㳲��N��褲X�����"Mh3&(6m�E`���S��j�o���܆x2�E���@"L|l�7T�"�)CkHTv�Gi9%'�1urס[����h�׺�t�=@���g���A��A��"�Z�˩�#���BEƌ?{��FEƿ�j�\������>�+�v1o#�_.�ʢQ\-�A��4-I��Y�%�����= H&�����Q_;,�O��*9�*!osk�f�:�:-�;����%G�L,��_���������;���x@�>�S������f���I!v0|�m��Ӛ��Txw�����P�������c[��<3���N3�d�N7�M����NT=,��d���>Mӟ���mԎ(x&�LX�d~Z�P�L����y�i���خ>K���]:���P�Z�gS�e5�Gf���i�3Ct �Z4���e��LVL��9/�:}��Q������th!����B�������D�ѯ�IW~���Vd��'y�����Nw��W)t�U��.�(�pl�ci��4'�ɯ���OS�ut( �f@�!Z�� c.����E܆� 9�ӛ�;3O��S �2e�;�?MK��`��a$,+���g��x��P[��ž���[f�эC��	L+`�f(�=�
K��g����c��/�:"C|�*���9}C���^�}I�w"�N����t��[DS Mw`�jy�!ʏ�w���O��4L�V#�p+t�u�%;|��Ą�������>��?�*�_�!50j������Pm�T^/@��4cN?%A�Oo��8FO������.tVK "W
�I���Չ�t}�pv	��Dt�����*T�0�!۠��@zdx�j�F(�5�b<��͘n���fywߌ� Y��e�о ���|�ͷ���.]I/��37�����مI�a+(�YL+i��)�U�Ӂ�u��xT��	6K���V�YƳ:G�l)���� C6-�4,L�>��1��5�y��X��e;�`+���҃�e����4�,��6d��K�tbl��>�ƽ+]�F�(m���Ʀ4�<=>�^?{�qYH�	 ^����9=��fdjm���ޕ�-
dg����0QAо"$@P��R4�Y��Kݐm���83(�p�`1B]���ۖa)?2S$�(Z���ז��G���(�&���e{e�hYKv����LHs�����Ҫd��U�F��<U4 �{�|�N&Zo$ ����n�L��2�s5�v�����9X�L{�q;�LD�1N��^��UF�� �h���$#K_� }���>�'\7����� ��fv^Z�T�z;4ñ��A���y�©w���F,�R�#����pAk�ֿ�yY��5��$Ç6v&|_�R�J��� yP��
ݐ�d9C�������=;��L�G)f)z}U�E��2�r�H����@���T	��g�k%�;;%t+���(G2��C���f�Lڵ���щ��v���]�A��!n�aZ#������ɴE 2X#����4��Y짘̗�n_x��0F�S�b��Q�r�x�6�	�pi>��K�̉�,��)�H��u����oa�>��ң�W(al��ޜ��Ȳ��R>����}4E����*;�u�{��y�r�T5��$;?��b�� V�l�V��������z̖>�o; ��o���1� jggq����X̺{�
�I��ġʱ�"̵�Pg�p$��Vz�x���Zzz��S���o&��w�6�}M	�w����M0Ox���+�4�I�i�"��e��~ذ=ڢW~��TN斔�$���y;]��+8H���\Ts�*)	pN���G��v�v藦o�X��цߓ�Dz�ѯ,����z ��g����ém�����\V��'RKkgz H6Y����.��PX}�E����m�j0\d�#�0G�,B/�;w3XlpϷ'��T�ǹU��խК�֠1'�����q���<�5<�5�����"��;dɰvǀ��Z��Εՠ�6(M������`Tg7����
��0K�xJmQ��ũ&��X�ݬTlG�wtE��u��q�OU���j�y�GU�$������S�t&�*�-0�ml2/��R���lbL��ݺ��Zҕ��n���]`q��3N�f+�ֆcϮ-AD��kg!´��gI�����!���Œ���F���|z��އN�}�a���&�PNè�r�,��� |����9n̢��t�����FQ�L��2��`ى��.0��j�v��3�0P6C���Pp�gQ}ʼ|T/	0?,�<k~r�I��X�2�Bĭ���k\�+ \e\sY�=D��뼈�|yE1���Ly���P]��0�z�l���ܴH9zny=bq� e�>B��w�J0����������sl�eӲ5"k��]�@�E8{슫=�l�����.�o�'�l���vaR�y~Γ�Wj�  �\� �,0�����y�$ �JG��w��ާ�{+����k����m��NU�vOK��ª~�	�.�hG�{�-<T����yX|x�51U<l�%��:A���C���dG���ω*�3��&��W���bUC{k-�g����f�I��]��#G���+9�����/�]t3�?����p1 ���_9�&^9v.�h��Q1Y9;0w;ýhV����g(����	�g��d�:K�|e3���4���
���N5�!\��J�9�ξ��J&K	�vi8ɱ.>��ϟ�n�C0J���E��@/�
j#/k��?K��$���(\��BٕvΝ��E����/����&����ʷ����F�l��啗�u�&����Q�[���Nyb�:W[tl���ܙJ�z�c���փ�h>���F�9Ρ01���g�ӝ�?�;M���ʩ�^�t�>�,`��a	�X�e-�����N��Y����R�8���!�����2��y�Ct�9�Ad��]λ 	_�˳�;К�uz���u��%��G�e��p�o"^�x�U��'�uƂ��rJI�,���m�TE��	����,���C`��g�w �,r���>�]ی�-������q�ӭ��k��=K�,�ӈ�����^�d��лt�T����`��x/M�lav�lЪ@��q�Р_���N0��+)�DL��O�^�F!��\<�$�����:.lw/옌��O�0P���SO g�^zeh��ش���A�2����XD�Ӏ�^���,+R���GK m��eIB�����v�1`����ࠝ�lW��v��,o��P���a�:�H5Tb_����?p�^�H3�l�8f�q�4�U�����c+X�����È�*��)6P\7 ��|�]d�����jԳ�n���d�F��n"D5ւAUx e��l$QK�ЇM�&�/�JA���wpz�q�W(��l凱܆ّ�Yۈe~d���h�x>Z��赴��O~�rm����+���fS)c=����ij�O�*�	0�ꄊ�����y){4�̯�=�lJC$��WY˼���l&��:ߴ�{���YA@�9�3�& pj0�+Kt�n��9�ԗ�:�O&b���z��#�n#h����ĸ��6��3�2���6�N1�K�өB$�dHc+.t�` e��`� u��
�ͯ�^V�I-������E��F{�Z�%��^���F}�D�}\;Y�*���5u���6��C�j<9���gC�e6a�5WE04l�������=D��6x_�"�[R���	M+�+�������Z�cϦ�'�b����T�dq�����~�C�X����:�2w�}B�7�L6�ڬ����E:�"��x�P�)�<����l�z��?I3\�I �F��x����CO��Bݏ���Z��_�VZ bc�JV�c�TPűL>P}�);�����KY�(�L5�9�4�ΰx��Kv�b}���n��������T��������01���&q��a�z0)�Q
i�M}`�yje�Y��p�rZ�\H+�b?~H�ߣ)~�7�]��vUh���ۨ�����Uh��e���B+�x�.j���c�]Ak���J~�������N@lu����}�E�����z,�"���A���
�ll�(u���Hc�����܋��2 *���\����`O�LJ]E�j1���Jt6.�2��HM���� �(�t�(���9�9Zߛ�S������H������10Wa�9r��J�����ǤϏ�[�����H�����3�)[�}�5w��v��t�έȨk$�S�̓*|�y�vK�0�ϐ>/�:(��eG����0Iu�[��hf��S����74�����(�uu��58��r\���R�]@'%E����JY;�Ԭgm�ټ���=:�XMg�R(1N��}�Ǿ�R_� D�0?���b�ǯ�	 Vkd�Z���6u�x��%(��d��H!]�uk� 2wr,ӈ��?@A�b�wncs�ᥥ�,�N��}	�xUj<'^:'K�YWk�y1�+�V�����V^'TAplGke:<؞���s��v2�!�)[n9f�\%��+ ���TR�+��jr |:Jwǖ��=��"Zb&B�+�?ňqMйZf,��	�u��gK�����k�(^���lF�0k�:׼\�M���z0��|^�k�=�Xc!1*^&�Ps�����3�dVA��-�F�M�D�d䃫����J�jkHsf�ٴ�[*x C ���Λ	����Ag[�g�ҍ��=k K�&�+�e��lA�B鄇�������L�OS;�v���t�5�I��ߛ�ם`j��6���|��;�=m��,�M���������n���!��, ��ۑ3�����p��(�	n��Ran@����=}O��W��"��G��mт�LΊb��J،C ���<�c��,�^}����������n@U�5����}\�ע�l���<�SbӀoƩ��\��\ׁ�C��8�E;� �b�x׮a�'�~7�O���3��y���ɂmRT���!��ǹ�����h�7"�Io��ct_MsL���K�0>wn?����aĽG�Q�c;_>WH��:��`��sv˒��?��O9�h�/K0���a�L+�t����s�2�`�����P-����T�pm`Y��%<���!3	�+\�u:�z)+�!�׬�(�"��~7�8i�������R�ևy϶Χj�R�g�Fpq1��˟ߺ�fd +mn ��y�����u)�Jm��;`��a�|V t����3[�'��s� �p=�|��g\u�դM=yf���k��� p�{��^�R�T�,�d���݀ylq� �2z]����c�`��더�,o�)����Q�S,n,FY]�i�%*��q��S�r��`�n��գ-����`�5��
~>�k�a��M���Qyemt�8ڟ�����7�ݫ�[�����V�!�0�����~d�@������hmɺ��.�h6a5kfo-�_�_�����EL��d-��qV�$WF{Q��j��dkv��[1�9z���v7��V��Vf̶;�i�"�-��t�L��f>+�����6������>��,�9VY�k9'o0��SE�n�,�;�ޙK/c[��ɑ4�V�Z����;����/1T��;;v"�L���.�a��5\��si����=�I���Z���ݦ�Vf`��i�Beq���4���rLI�XI�F�X�*��6 ��ڀ0uB��Q�����'ЄuR���Z�U��M�_��/ �Q��J+��ؕDZ��l����Tg�#Q�#e����r��4�*�5��>E5��*c2(��>'�; �<�P�+t��̉��?����2�t�����=�����3=�c~�2��[z��A�NK��&v:mB�m�f��x-�YY+����D�t��:��(T)�c�w�����Q�������,ˣώ]O}���Q��R�h�M������.<��̖z�G_{P�YЎ\8M�=4h@r���9�������oT*�n~|2��3��� X�DyE���'	�T��ț��sv�m���D��	J2���i0�D���B��E���P���,��{�l�{�N�G��/�ԬR�`���<@���O~נ�R�LQ7��$��r��8���1�������K<���q">�)m�@�\�6�K�^IOF�踡�I�	�P�M5��;���[:������n؈��a�b��M�h[�(���/�9�=c4[-�G����2�k`z�Lfb��o}7��g�.�>%��0�l`�k�Y����~�FIE����2�� �c�;��:�{���\�Xl	o�)�e�?��侍�x����P��
��� �^���o��Mi�����Gt����SiY��v+�[�}=����)�k�>��v������"�ytW3������橀�b�]s����I]�������.�</���`(b���)��P.�1��/������ִ��i����E�q����'˱���n�1ҦIW0��`mid
(i�޹�jas�af��r��dxo���3ҩC��)]b�D$��Y����q��Ϛ/n�h(+f��m�U�෸Cɚ�Y��<���;v���%���#��(����CFIƁ��m��F��#�ъ�Y�w*)�-f�@e�Z�6.�|-2,�i`^���Q`4�;��u0��h|�����R4@�r���_�.3Q�t�y���@��q��P��)I�͇:�`+��2��e�d��7r �r�������4���v>�Zj����f�(��L���v��&�j9��P���d �+�#���G�3�6B��V"�G��JU�NՉ�j�ES��f��T	��H~��4���__�x.@��T3�����_�����K�;At�o�3;p"e�څR�Ci"�b�vL)�����ꐺπ��+պ�E�	NzY�u�R��%�d1��� k�����IW��#�����.ϴ��]-v�1����A��"3w��r�t2�3�k��,�p����	)�P���6I�/���vu��0��Y�E� ;N�v��ٖ�Z1'<���z�f�lK�YpR��X�^H���I|~
��ΰ	֚�r�� :@�4���|�<�	'�
��aܑ���ݻv+]e�p�]*�+Rv�kj1<�f�݇A�F~����:�cZ�7p��\�/Z��r����Z�YTg����˲�&i P��N�M���f�&t�,���[���l����0��CSV��0���u���A�O7:��ɧ�B�yE	�`������"����?j�k�'��s?�B-�o�d�pX�$jce����(�Bt�{�cZ�g�-�R�,��uf�J��� �;�ǱA���F^s
v�X�"\[P�,�E�G7�ћ݈I�*��j������ه�)Ǝ+O�F��5�S��s�]���+�`��ǽ�Ðq�C�� }%���b����y�"�]��%���azG��1d�|Y �
�C��x(���������1��k�h]p6 �������$�v����3 �# R$��kj	��8fm���9�Ϗ����f}�vz�X�Ky�}ک���C�%��$���H��J[��ͅn��6̽o�91��%Lw\���:��Z�o�a�k`	��d���UvK&����D-8v��o�IYi)��3'dE����T�_b{�����O1�:D�I�\?��Y��?S؊�M��;�3a�m������i6o���4'0�$Q�����
�%*���A������A�@��I���b\Ur��"�� V�>Jb�o��6���'[��2wt ��&�0�4Z U��2NX`�����)*x���?;I53��q�ʦvҜ�����X�$�y������)�X�&���<L��ܫX�;����x��zXr�ì05 #���e�0Z����:��*f �����M��_��/ �Q�r�>{�x$py����5�Y���L��Q^��5`wa$43E�⥌���v)�-ih�������!��A�U��؁:�`Qt�����z/�]&d���b7��V�M��w��	��zQ�g�R�Sli�����^�(5R��n��hfQ{�嗃����Dh	�߰M��%}K'ݢa�zY�uB�a���믠�!ϊ���b����[��X�&�'�Zy���'ij�1mĳѽ�r�S����= w]�4�ziy!�6�V:����4�W�dQ4���{4[<��t?@���iG�������O��EZMS$�?xp�Ũ��o�U�ٳ`�"V������4 N�5�g1�<s��V�'�cVV��|��|�I0;- �]@�e��@\U�tm�H��`5�yZKps�45��=���ьP2���X���>#"b05u��ԡAaW(M?C��&���?�#�Y��&m���n�-�}�)�-kBi�?�d�]:Ϊ:�L�`��� B[��S��D�0�7�2ô�{����IJt���
����]n?������$�J�@�Au���G�n�ӗ�"R�>�pih�ptCV�SItR�D�L���p!\�\�T��t���0�l*��`��x43wfp������O��R�"��8�Ȏ<Z�ZM9.�L�>
�Qzx�����є�F�q^C��`��M�92�&�'͛+�N(�X_Y �Xk
[�ehؼX	���*�yмs��<]cl���d��4�S#dZ}�R�!ȵ0��.����~L?]L���X��o|�~4.�.�jHR}2�r��q:BQ����u"i�Zr�_�}e�[rł*�d 4�f�h���\�e�ik����@��ç���3){#�	}�A��s���Q�	��ټ��ZޘB���o���N���?+��51$��-%�졛3��s�H�'�V������p�!~"d (@׿��Y����
�����tU��yb\lqo�^ۀ�9�66y��;� D[�Ȣ[B+%�ÎT=�.�-�w�������^��,[�3�M��F�ȿe 
�M�;�bH��0!���	��3o��G�O'm�q_����s�b�pra�Ig�����AՅ7���@�[�W=-���c��o6Ѻ�6=�����&u���}�=����Ձb�ׇ�����MBC�dj#`��,M�Jy/M�|������Y���	�	�H��s���v��aLX��-B砐����!��������r�� Nb0��w�I�#�{��lݒ�&j7^���S�PبO�;�yڛ��Rҷ��.vl	�$�cvxL�Ɠ	:����h�N'�x1�޽]H��Z/���dfy���Y47��ܤ��ݗQ2X=q+::����!��t-���
cQ��+�=H��!��+���6�j�+���(�}�jA/R��ʵ֧���4�����=�G�N߈cq��럓��������X�F���{Sc�Yj]���iܭ���}�R��,���u��)�)�(5O���t����)���y���4ȮYFOvd�n�y@ќ��k���h5���HS�Ӈ��?��"���AJ{g^5��� ��i����.}��n�̏>�[��d�e U}Y�ͯ���?x;5��VCvq��I�YP�CG��Y�������/~����(W�*����!��n�H�>��Z8]Z�,m�X�[�����?H=0B��Q��jhjFp������x�R�Τn�|V�C�NK��鵜�U���X�'�[������V�
��ĵ���o�Z�ҫ�S���<��\����$��=r���	P�"g�������������Z'e�����[�����b!e��a왡�g�b�x�u}_D�b:s(s[�}���Q��9Ư����E:?�FS0��Ռ岥�Q0�&~͂��"۔�me�@��u�4�����^��n�e�}�N���<�l�p�����Ȭc�I�Bdm��:�P#��E,Ζ�����W)��˔͙�=u+^'�ݎò������`S)r�}e{X���T�� ^I1��A�"}�&e 8V�4�tg�}�)j@��܀����	����L3�s�,��I6�%�j��6�C�I�;�	56eK�#�}M5n��D-�C@

 �y[��f���cQ��u*;b��rg`7��HFi�.{�	_D���.]m:[G=�C��.���5�$���}����: �#��`�D7�Lֹ3:�	B��I����t&���.D���? ���6�e����G�l��?	�����h��ά�a�RN/�@=� � �T1�y�G|����h������n�yh����")|�
c�AL��!��(��`����K��.�~"kޟ��>���ν�� "䩙�(O�q��D0����e��[g���4W��5��d�.iM��׮�G��H�&?_���Z�ڪ�t�2�G(8�v"�9s����t���t���E��	^�y�F+�9�v���d,��_�;6+O`�%���K�҇�u?���cgف�L��ꏟ=��1;�u�]ܫ0?��KD,j��&g�����۩��l�%�؉)��L�ogy�����)c���12Ў���]:�`���_�|D�����/NJ:]b�A׸E���-�u���Tz��4KԌ�)�P�}�� �S�M�����v"�~u�i*ÐqV�����C��6����ɼ`Ss�����1%��3��O���-�*u�l㵅�ؿ�7��
%���.B���k:�f�.�~�S�\���]�P���^D@��b�Ә��z���G����a��u�J�l}�q.��~5r���?Lkl0,A� �(kC#6 �墻N��$^S�|�i���Y��:KiU݆����z:s<Z�� =w�}��:h����6�ܚq����̸���Ȩm3����B��/�8�j�W>�<!׭�{���v~���3��7��a@�*�e���W�5j��8��m �-ئ-ة
�GC��:�Kx���(��o,"��yb��P_+�n-��w�2H(W������M<��`�\�]���L���N����\��NQ�l���g��j��ԙ�2���]_l��`J�n�����v�y�#{��)6�� ���fT�]����5�>��e��\k�f�֡Q���U4�K�A��A_��.��5�P;t�}�]���2}e�N�=S����0�:����|���6�p�M`P�l���a�3̸W��� t�v��ls#�|���iI [
�v,�gd�8w����r��]`������n��SOtP�uA��؞��̕�lf��P�Yn���W7`ؗ���+� /ip�Q�=����eƉr�z Z��`?�i t������,Dp�ё��.+S���Ο�k<�~[L�L>
�`6��ja�X�,��<�	C=��fv�Ͱ):�u���ؽ����U��:��L�o�1�:jK��I���]Ut��ðe|Q���5 Kһ�6鴲C�����,�����������N?Ay�Eh�����7G�����f�b��\��,�N��0_-��#�.C��;�����v,��AJ7�L�*��YG��Xc+e��,��쑵�|�pj9M7�!��K µt�(�E0E"�ֶ�*Ƌ�\�9�a��׼$,l��-�Fm�8�;�N�@��5܉�(��G��$%����=$��^J�]��i"��#����G�mHKud7�iy�Π9�O��o�R�����B�;ۥ˟�q�IE}��}���[��������C8i�v������W_�8ʲ;�̪�9�����t���4�P;�DI��S��* �-0hU�r{����i��!��~\�Zv�U�Y��;'Rn~:D�����qv���=� ��l;B��*���F;�z��۫�l�K��4�������mm㌡����͔���o�����J����ZZ��O^|!r�0��x>�(���\��M�*�aL���/�M��3Q��������E9r����	ygk��:���k�B�3R�sS`1��1���]FL@���X1�_�a;��5lVV��G���t0J.pj�X�B�"[;%<�(�L�f�+���N�q�`�r����� �嶉_���_��T�ȩM����i�  ��y��<��`B���,ӗ���H(S[W5�/�]ղ(�<�x��ϭ��Ñ��̔��N0���V�J��v
�*s��s�KsόΈVxe�,�q���KrKhS�Q�=���?�{G��&�k+��9��WԸ��%���xd�-')'xZ�P����͡y�d����`�\UCT.̻lr�#¢���@�H��>�'��|��C�*+I>�P�fx�J*�q|ehA�A�>(��7��� ���e�QD�j9��;�c~ِ�վ��E^��IFV�Tظ�.>�w��J��(gGU���m�E���*l�����>�v�(5`B�Eo�"�[�oo���}k�*��
l�����j�.&�>����UO��\�6b&b=Pt�5����y�n�+�*`��4��c�$�v��v�P��ֺXBi�	�B����way.����}v=�O��'#�xS�]�z�� ����ݭ��l�P-!�Ns�WS:��1&@J<]ͩ���=G_l�\���\Vx�q��L\9&��0.���!P��%�����[�� &e5�a���:)+uVק�~�^���Uf���N:��)��n�j�,��oR~:IًE�<-c`�i�& ri+�ÉXv����U�k�p�e�p��2��;D)�m�<3�e���F�_D|\}��Y�`�������JM����D�3w�jj�~�]�s}�V^D�5OX���jF`}����`��b=i�� @f��	��LQ��&��*���u8U�,��S�(h�L6��c���O��s���9J.� �f�s����v%�nW��_�}�na�� [�C�"��"�&�cv���J�ο'Sԭ����3�	���]>����fL�Æ�c�I�����:tV�\�}>��7��E�b, s�a�ƛ�u���߻N��~:u�Z�%JP���9�Z��D$�ä�)دK��T��:,(Z�.2�ڹN��� Y[Kt~1�[#w��A7zA^,���׈Ҡ�WO��œ��?�O�ޝ� ��W��`]���VЁ���� �L;/U�.&@��ܻF@�ڠ��.�Q� ���NL�}䩲QPl�+؁<|_o�8�V�+%���#��ۀ��0T��`��o��r��1bێ+����&4Z]ca^u����,���5V8�K5hD^�b����(�g�Z��0݄��gN����g���:gM�"u���$
@��G�2.9�f	=dK�,��s�"y��J����%�U���,2XA�!5�^� $(A�T����g1�2�e9�#[��0Vel�%-a�+È��0
;���S,cf��k�g��U���*�\��R�[.Z�? �6��lqx.f�n����c������5�C��2��V�띹�XN�<̊S
�l���)�>+� �M���8����9���%fʁF dwPUAA!	8����d7�pv9�ߜ��2�����N$Lz&�����p�\D'���k;��%L>�,��<$�'����Hy��1��H������N ���k��p(�W�� �6}���Pm���g��HG�O��\�)��i�`�.�]BF���`�7�v���1��q"*fY Wimv��c����D�Y3L���	��g�C���.[��z�:f��)�v=�(p��c"(�@KW�3���-d��#tb$:ET� ��̟B|:I+��̵�V���H7)�"��qn �chKԐ�����������MSʊO?M�o�F`����&��9��A�}�JnPk¨�U�L�cA� �R̹�gӕ�>��ݥ�t���
״��v�j�����ڞ���/|-ė�,̥�����������4i�~��!d��̭'ib�a��ӪPx
`�( ������:K.��ػ�ͤ!��\������E���P���h�/�?�w���eg�������2�wL/��-�W��s�������oc�Z[��ۏ�(ׯ���?HW���n[��ǘy.2������Ɵ�2��V*�Z���RloL@������yV�8�,A%���A�Kg^�@��#M�����E	o���1,���#�+o��݄y7,〗�f7%0�aݔ�ԝM��u���(m��.f�'�T��-W4���l����<�x�|�D,f�0au��T�xml�2�HL@��,X̹��t�m2>7���sj��dq>��)A��N�8��S��+��ߑx���֢D(�[>�,#X�D\ђe/5������}\��{���\Ф�ؾ�^��`Mr����R��A� ������5�.�Ne26�
r�ԯx,e�3�g���*�/�üTm�Y:�I�=��ĥ��!��=�gl�bK^��g )��7 �nq-�xT�=���'�O�2b���VLf��8I �2V�h�v LE��m��<�Г�9��v�uƷt�u.��HyW_$o�Z(���aI�B��6Fi�p�4CM �M�zL��T���U]t��@G�+�u��]i�Q?j ���Ysv(�)�gs-���*���|q'�\� �:u�[Qgg�G/B<�j�Q�ˠ0�� �#��`�[GHW�=X���D��ԙ��pkh�J�8�M,B�+���Z��Tm;��}�i}H+�J.D��i����F��A��s�F����T�ٴW4��D�TR�Q��������Z�2��jX�K���ޢ�0���W�i ��@Չ�k0`�eZxO_�H��,
�i�]�vh$��4UԘ���+L.[a�7E���?N���(i�Tlw��S3L,�:�Z�^�&�F&1���N�=�ߟී�������MK|	�����ʷ� �A]�-h�f��"�t�ܶ�$��Q��)Bf��z n�n�{05���~���7���4������	�����$�D�����SJ���m�1�l�li'P�F�,�/~�t�������l� E���w�.�O��5gMWzB����M%��`g�>A���ӄ\6t`7p5s�e2~�	�0���������Ǘ>��`M��G^�Z}�(�g�X@�0�+'������3�CG4�0~=���ə�p� Z��(3������./ؕ+_�](OC�AT� �g)��b��/�>-�0_�Zz�O�<r�,UT�d���+�����fqǳ��6���[���r}���ʁ=�fگ	ݼ�N0>�����`���,ޕ�?�!!�#��{��14dm������EL��k�㲃���X�[���j�tA_b���5F�c��l�l>��aJ��o����cbM^ �%ǳ� �X�� ����8����R�����-JU<����~�ҥTa���YB9�p��1�g::a�:(%ʀl���2��v�������h4��ǳ�Ƈ2P�f�+�"�<�p0�,����虹��A@��T��wKK��R��N**����qa.����"�`*�#5F���s֗�T�; \�j�
�:cNz� �x�g;zp  =�,�	��J��hW�$`�� � �<�at[E�s�*�0+�0_�[�`{c,���m�� (���`�'c�a5���I$ȕ��t !�}�{f��>�*U !7�j�L����F9��uY~&�62[;�PX� J�ȪEt���ʟ�<���3d;�6ǥ�A	�dPQp'S5�e_��"��s��<CW�ٓ��Z�}���؁��}*w9{fr��5ˢ�P]�������e�]o�;�t����;��bm�!�T����2�N��Mv���Ќ-�lr0sh�V�7ݛm�uG���f�ؖ����tF6��@	��O���b� Zʻ
�N5�@�u��$)�AJAv�4�s�6�j ��.�5��nV|KY��{����/JY�s��>2�-ñ��Ӄf�!%�I��m^��O7�}�6n�g�(� P��tF �M��.�6߲��޿��~�׎#L ���o�?��E�]G=e�f'|��_�j�DL<���> �T��ѽ8o��i�ڍ�� ���J�0��������jdZ)C]\�*�����N�ck�ª��4{�q�ÄU���b�O+}e�:b6��� ���@9�(m����9����T����Tت�l'��bT
�Za��$�j����T%�d�Ϊ>�c�'}�7�*�x��0N�E�4��Ǆ�dj���Ť�{� r�ֶqL��ɢ7�d����mP�5��v)t�q�q����T^܈h�etne[ӰF���Q@^�`�tS���c���B+��c ]�+6Pgw�I#��[��� 	��$��g��w��x�h����b��hG;Z,O�qc�����5��1HT��~m�NF���Ԇ�.Б����1Ս����I��j8�A�Y5���F3ꞹ����ŧ������;�y��I�_%�D���+ȞrAS�j�CM}��=�Yn�Y� ^K���V(�k��|���DO$��V[�Ku�81��܃v����x�EJy�	�-ߙ
0Y�X��`U�\��������cU��q�@3�D���EٯJnF)8�
�\������sG��dj��6 �Y�[*z�L���:�l�Cl��s,B�M�"�-+��b�Ni�j��%2��o�d)*�UҤ�}�A��!�0oK ����b�:����Y�@	�*�g�U��k<k�ey�eh)��@`�(sE��j5�x J�6�vl	bD;e �
��}�����3�-�Dڌp�"�(J�N�R�י���c0nF�,+ Y0T�2i|�csMȜ����\f�*_��®�s�q��Y1Β�}��]��١튚�*��s@*�Π-A���){X_G�agE3^-"�Zk�v�Uhj N�>�%h����<���6h�@�L�ާ���8����A�a������a<���̶n��Ĵ��m�N�Pp�nK� d7���s��4����0���x8?s�r
�\����a,+4��2��Ѥ�X�J>��7�Hmh;� ��w�h�ň�	"�>Z����24���s���'��hA����)i�e�-hƸVҚ^"z�8��%�V�Saq��|�� ��@_eR=e��~�4t.#����&�[c�i�`��s�Qۀ��чi�����Pz���n��R3�w.ޯ}������,����ȩ�MGz����M��3q�R���Q|qZ��� a4?��\j�us?�>9y4�;���`��b]3aP�`�
���� Z�fa�^�p``��b�w1�&�c8�܋V�v;��E��O�J�����z'ݿ|�l.ݥt�xx��9��M&�܏ou^�,��y44�����`-9k�S�W����!�,��8Y��A��I'��|7���C2�zf�>�p�ћ�M���b������p����
PW�,�a �b������ ��{��+]�s�Z��9�Z�\+�0��H�o7�0p�.�������1|��46k�GYx��������U3&u2��% �)�]��BH͗��E.~�yw��,U�k'�[����p(;�\Â� ܚ��8ЩF)$q��@���뼏�]sS. ������5���b�kB �f'���Yh���څA�<�	;�\t�~��Ȓ0�M=��f�K������߽
�ݱ�˴7ռ���ھz�(,5E�� �(���l8(Rt��r�vHS!.bU&����
q �
;���Dk��i �g��C�{;��Nu����a�lϚ�~֎2�'��d-�����ڣÍy��U�I{f|�T�5.�X�
`�F�Y��m�*��H�j�ST� ���JOs���d��G i��n�Q͎�/�0���GΤg���{!��{�>������������E ���q%�lJ���Ŧ/l����
< �S
=�-���;*�Q7/a7�o�%�����0��N�yQw�Y�K���k)�UQ�X�m9���i�G��G��VP�n�[�OuqqR��ct'u�N�ȇ]*��D���.�զ���8!����LU�nu�1��+0�����t������g�h���ٳ��1؜bx|ئZ
ſ�{m�(�����0����|��8m�\�2���NW��Pô4�(4t��*4����ݺ�S3��,qlSʸG9j��v�]��ob�w����e@��,�-kLlM�;�������zs�sWG�B�kb��_ݴ{W����r�|�ޙY�x��tV]��wY�?��]�q��4u�n1X�
���VУ/¢��\��j�M�_���j���@ۣ6g���YԶS=�]��R���h!��To��;�<����c��6^L�.,Q.�]֔�;���Q/1��5&����"b�[�D-'��؎v�@l9N���》��ަ�ގ�����ݴθz
X����O�WLf�k1r$Dݫ�kw�͔>��KX,���_�����WS2<D)���wn\N?z��t��R58c�����+_�J��|��oM�y�A"|��晹(�X	 JY�O���Dy�h����g�
s��+���c���c;�}�˿ńsu=��t����µ}�x��g��q�^G�=�� ����Ov�������R-^�����믾LW�ٸ~�w]��CX�O9��%va��Q��
bQ.��!�ԇfj�<7�[�Ο���H�b--���5͡��� ;p��u����q�&��t �bF>X�M<�j��PD�� &EJ��&�h�	ʎ�k�nE�R���>;���r���\[��MO��\� ]�gČ��C�k���ܓ��3��H���)5���V��3�gtJ�����yU&�?�������Q%,������s'�C�K��)�`��MW� c������0"��4�M�r	c̬�L���M�Z��(?�����F �G��3ǽA�;�%�e�v1oo�0bѕ�9�����Մ{�P��wYk7�v�1?��f��z� 9�\�J6�:iW��yĵ.f`�o��w�ԍd���/�
</ HZ�R-R��"k�@"+������vaH;������D�Rb%�y 
��p`J��NX� �1�&��5W�-��Fd0)w�d4��;&'�-v�ch=�WՅ���n�6T����w�]b�`tR��;��C��١�k�>��|�K��f~]L��t���,c�]���j��" ��������o|���� �aZ�#���ha�߾M��S�z<Y[,4jS����:x%�������Ѯ�@��@��mr�rxt�y�sW�:	��z�0	6QR����E������ǔ��q~�޶j�f���}�n��?+X��9Ƴ��5z�Y�������IEyWZ�%$��}��0s�f�L�%|��_�aU��PC�M$��f�,��481e�����)ƍOFoB�/㻳��L=���/�љU�k�·(�B����Bl{��U�1GB�9�?<N5������cxlw��[�M��u��%�a�v��sʵ�`ua�G7]7%˜�G@��9�B7S�=�%�.�q[t0=x�4�Ie�\3�R����/� KF.�~�E��y�.�����wñ�B1'�|�����Z{弭2�|f5�¤4��|�si��ߦ���*�E˻��Z��s�&B�5Ev�ë7�mX��J��C�ܖ`���,��O9�6q���֣u:{�;cu��Y�st�֭ȟ;5r,P���� �a�i�o),���A�>Fh<K9�p���K�S�g�Kh��u�-�$��1(M�n���+l��_����{��]p�%leC@�I�	�:���R�l����0��9��<%GJ�</�pH��+�Ҋg;#N����!�F�s�)e��>/���G��.��r�gK?k�g��>�Q�/:�ʂ�r����Țw�Mރ�+����{m=��ć�g
�p�����m�g�;����0Gd��Rf܄_0�9e���KoY����9C���̳�^����s�5�8z �����(���e6��xXf���f��s3[���@*aiݰYlH�l�#i���810�u:Qd��*�U��_����xQ���,�i�"	��R\k�C��z���A��#�n�w�zqn}	�t�K��˪Y��@Ϳ�?���2��H1��ɇEN.�lp�����J���|���P��7Ǜ���{��Z�×9率�C�{.@��&:C��Yآ�]�B�/bw�d�q<�5�����?���� ��vڥ͜]q)�G0�m���"0T�v|�&�>�"w�A3�&YD� �b�;Ryp}Pd\ܥ�3�>�	f�g`m��G���i�:���A�Lk��c'�|��vg��a��YD:Y-�5���]���]tp��0�i#�d6|^��YkPw�R�ڧ1ZN a!z(��2C�F]�>��(e�Gw؝s���t|��/���j�|��;U�n��oGZ'浵jR�����)Y�౲���]��鋩�	���;k6��h�Ώ����i@�N9e�re8j�PT��)�jv��#5�^x9���k��mE��ct^�6_�<A[��P��k�NQ�"n��fX�rĿ�,���x�c���F��t����hA�+cw�3���ՙ�g����|���S�O-�[ GjQN�
��9�*���\;��3�qo���33i�RJj�tB-!p/9���?�r��!�F=0$�m�=-�M�x�ƦR/�t% � �����4�~� ��>�8M߾E)����Ck/�ŪM-Տ�	e���f���&�[��*/��`!�)/�s�Pk���4ci1��ߧ(;�n��4yf���pm+�Ǣ'��Y�-��[0^:9k��P�g�Q�5��݆)jB�eF���c�?���YK��2A|���1T�n�*�KQ\O��]4of�	�d%4����..f��U�t���Y�KH�?��	������tW~�(!��(�C)�#@�NƵ,��x�5�^d�& Z��2��g�'�mdз'+�eF��#��f�� ��a=�t{�,��|�i!,��,o��j��L4T�[����ιEߝ���Ɇe�^��%.b�Q�j��dZ,�d��h�J�-ةh��X���6��Q!���9�#zP�K����9���M����4�0����v�RL��9�:���ճ�^�i;�8>���[�����  Ja�l���\U��N�G��Z+&oKm�񥉤N��*q���֋��.Ҳ'���8�9��E��r���{ʶ	&��{� X��ݝ!j'wv�F���k��Ͳ��nE���g���5.p ]@�>�&x%g�0�!ش�!���7���ؑ$�XV&8�p[�+)���q��޽{wn����O������z.@P�1�锖������s ��
[�8b�DY6�w3Y�i����T|;< �XY��9�Av���ԭt���&l5L���l�fGoǁ~#n ����C�5f��u,��*K�I���k�j�M���!�v��l�	���������v���:�*j3���L�����jة��E��S��J� +�v}g��s� %BKs�q�2jK�8�AĨ�#���ɥ�ѩ��;J�y���#J[�w���i�D�G������Q��J3,B'�C�H��`�������^:��H}FY�Y 6x�4�R��X��=�ȋ�쟥�+���:Ow�$Q �f D��_�g���4��8ǟ�I�K� ~2jC8��ΤeX�EX�j<���V?�t92�>��GWI� �p�;(��:E�ඌ~S@J;��H��%�w���dz��?�� ��"����s�]2��n����@� �=�k��%��춠�a֮��p���P����=�Û����{/uӅ�d6	��<}� �5�'S�'`�6�&���_�J~c���Y4^Ôٺn[�\\��}���M��)����U���֘~v�:��`�6h)�COq��_KmǇ��X  ���)]�󘉽:}���~?��iC�65���,��LЇ�T<ްIL�ͮ��薎�:i���y �U4@wI�/�n=l�����j�c��a��[_o3��é����	픶���8>Y �x�t���`���|���~�$����9`��-^��������A����_�⹭f�4QZ�𳜟�ټ�{i��WٲHdmB�TRU��csPY�� �X�)P�ei�g�[���aAU�R��Ac&,>��{f���)�u>ɴ@���S�^l�},�\��6��T��W���s��,�K���.*Sl(,�Ph`�ϱ���+��s��Ȳ�Ɓ[~��x���\�i�,��Ȳ�׎�MA�s��%6�YA����kL��Q ��C	�MU��
�9�̈0��F��9���F����*6��lh-])^���h�:E����4-�X F�{@��@c���<�0�����a|6s��Bֱm�R0v�e���ރ�ɼ�b3ic�`G�yf"�7�Բ�
�����]KK���:,��ga���| ��3������'ˁ�l2Q�J��YYM24V|�������|�	+)��ޣ����Ɔ���[����	��z.@�w��0PP�v�n����^�4�Y�̚(�~�3�J�6����<��0:{�{�\�D��n;Az?��`iذpn�KGZ)�P����x��EwH����9`Kaq�\Pl��DPo��� 2M% �8�1w����V(��݌�Q�v��>OvN%�h���"����T�������'쐗�$cY�����8�\�,�Kق�_`w>���aږ� ��b
������:ت6�叐�A���v�X�;�� x�9��f�tq��ԛ��`>H�;���	8fs��i5���o��:ʄ���E��jY�ډ�h'ꡔ]z��3��� %��ԁh��<���g�{l6WЫ<��׍e	�$�e*�0r��R�Qܰ��'��e�%�䘺��]-~v�-�ι&���\���I`�s����`&Q  ���t��^�5�vdJ=t�PF�C�|���M�i�@^ǝ��� �5i����}�F�(���W.޳ܳ�7�Y4��9 ��S�ބ!ۅ��ݦ-�$�u�_����b�i�� ��7�$(�8���;�fѮmV6����t���Sg	�W�� �Sj��4�Bٮ�,d�ѩVhC�EGڭ_�:}|���s�����i�� ��}����3~��Π���6��M'� x����s�t�>�lV�bk����Xz�������Jzt�z��·i���.ZԱ`O=g����~��r��C�v��:�!K��|�2�{p�����0ka�:�f���ѻqa�X��Z�h�a���y�e=hZvr�-Gg�Xem����[\ס��8�:���W��kL�1���X���t�e۪�y�U^�=Y#?S*� ���EXS��!�"7q|�'����-�n��U�˖�yM5�����((��Y�<��Ƨ�c���
6��"����h�d���-|i,��yF�T������+,�x�em0	�q)�=�cAU9]�2ҡer>�$��
p��Y�������,sh����2��R(b'�N��E@	p�����6�ǵl`���8ߺ�o�,n)�ήeَl9��=����^�R2��h0�e�9�Z~>��6��>��R�χ���x_9oi���W�W��d���ʶǭ\��{��)�V��*�Lm��c+��I��T�~~o�hd�jԭ[%�yk�;_�:b)5��F��(׹�q\���GO�,�!�3��PY
��ewib�Tf��{6����ױ�/�u5}	�~P ��>- Q����
���zz$�����ui�Gh�j�e���6���@E��>�l[3g'��c�T]���J#[����n��e��uں��R_�X~�_�D�i\l�EGA;f�`�6��#�0�r�� f�D+�MՃ�&{|�A~�Ha��ױY[�ϓ�>JG�J��^~�΍�S����ÇO��[r��t��x� ���z97pμ){d<c�ui�-�6��x�γ��E��zv��C>�&���m� ��S's�1�S牣 /ຽ0�[�lܼ����ZF�yr/�}�����o��iZ������|��!���xo�S�D�It篾�j�8��>�v����X(�(����/c1�����-RV��ŇhYJ�(k%4;�	A� &�>W������n�蛚4��r�+���T�I�'�:��+�~��w/�|�-�b?��/(�������=g�7�*��wp�^�A]ɹ/ �%�X����z�Q w}��*z2v�+0��0nE@�(�3KS�֍�i쓣0& ���]몓:@�(�R��E���_�Jz�1T�������r�g_:��~��|�`����-bT�١�u�8���
�DGW'��.�Ki�o��#ʟۜ�C�nq̦ ��[�{�|�\*2��身��Oi�zM��K��`-�(��aw�Gil �B��;���ۈJ��9��|XS���_��%lv����V'w���t
�L�W[�2�wɚ��уU������i�;����-<�d�� ���C��-����r��87<��#g^����Y�%/��='O���!���I�ߏ[3۲X�edHd��]f[�_��<�)dt�w��Y&��U�z�KX�NMqp��ZX��:��v;Y,s�5�S�?%4c*�x�#E^�� (<,0�e|y=-症��Ś�	1pV
�x��脝��2#����|���e�fw�-�%�˫eT�����m(�m�YķY�͆3����$��9�X�a�����e��a����%;�drJ)�3.4��ϱ�x]l�(f�_v��F��a	���Y ehr\/A2c��5C��e5�se.�6v�q>[TY)Jy�㖺�~�Q�Wqo�5k���yb�*��{���`mr9(����<��J"TK�4�&���e:,�L��Exd]��iR
��2�����;����e�����A��b} @�(30���?΄]L��K�H�a�4Ɋ =~d��X&X�㭱G���}���,Q-�[�X2ؤr�PGx;NK�
h���CE���>@�9�h�l��WRp�[2�u� U�3>���mL^�T�c���ux����@;����2:,�C,@��+l���a�<�8<q$Z����G�?����ƭ��g���Qh l}�2��N%�y����~�N*�L
�^�^O���~;�m����VX�6�0�v��$|�[�Is�^.��Ρ���y��̬
ص˴��cq7x�V{3�:`�Ыaa暈�@�r�i��Mvb{�~������o�j0P�F2	.�]Cx����C���[S��v@�������<Ү�`�^ƀ�{ii���:�}�N�d&[?����1ᖣ�*��11ϳx��>m�Zw�tQm�ץ��7�ܣ{i��=��������|�����"��� Q�.�O�,p�,�m\��I���l_�݄-��/Ӯ?	����d�L_2*�n���%U�Z;�Aˇ ����cg�s�(e~�"h4\U��X&��#Çp�G��n���(kNtU�X�E0lW}�%=��5���&�a�r�#@\gL�	E,;�h���[��Q�!��)/67����E��MU���@g���H�������z�����ױb�]�x����	�;q!���K��!�Ǯ��l�,�����"�=d�i��e739@i�-�oz-�m	����_�<KeL.5��r���fGjxH,���j=b��!��B�x���8+��oEw���3u������k
h�6y�2��
M]l�aU�� ���n'���Z	l����yǩ����7�!����=lG�yK�*S@B1�:ǕXVP���r��� t���d�I��v�(A�U���43T�@�<�
�?���,K��-o
"Lx�-/����#���!�i�`���Q. 2,��q��,��c��i�س,�n4@υ9�M�Q6��6�� �Z���@�2&L�d�lB������*W3u�	g��c���1J���Y`�{ܾ.:��r �F E�Hã��#4BY��^�~���0XW@htF&�!��w'.�G~�+��J�ܦ���|�IS���p��΢��{.@� {O�Ɖ':�Ů$�²���o�ʟ��ݿ;p����cHA���&���r�8��>�UK�C;e-��!���E��e���|�A���G�X=����lC�e���[��J�ݡ*#�	'w�s�)I�h�Gq2N\`�8�)W��"~=S����B�H^�󖥪I"��Ց������L�&��O>����l,�]��Ȅw&�ɝ��㈅'nߍ���ܙ�G �l���yQ������Ѿ4p�(��t[�f��t�r�*;xv�R��hn��5:�ڎ�H����M]o��ᐹ��n��6���{WkAحߑa�թ���.��p`>AvU��_���1c��(I���w�&��"Z��٥t��O���@C%U5צ��N:�����Z�+�-\M`�J����E_'����'�뺃����L:�Q7r.������^H}h��(�4��DsL�9�y�q� L3c�ivA6�|��D���0)�v4D&�[
:Ƶ��+~ǋg�lw��u�[Gϧ�v��HS�Ty(��?��R��K�l���;:��G����ޛ� ��A�B�]d,�,=}"m�z2����^>[�5^��?Ng9/��{����ϐo&�]Y�q�a��2ݗO26���W��M߾�>1ӌ����Oю�Ãz��y���(��g�=�����0�P�
�����Y>��l (|����`/,�/���j��ٚ#���F�,憥Z"kh�\��.���N6*��@�8���� �C�Y--����m�s�=�lf��5�Ayqr�ͅ��X���X��2T�<�c��\$@�ʅ0�x������&�Y���Q� S�FYo���	kj�Ė��fw������9y[@j��,�e�m�EԖ�xm5c;X6��V�%��s�k>�J��n�d��/�n1��������Z[Uk� J@#��F/+�X��[O�R�u������$�LMiy�J�s�� [䝿ip�	�������昼N���q�X�	��[�����c�k����t�kV0\�r��d�e�Ŀ[������iᚆe����Mg���<�9[�3��|���JEe���57�v��dG���,�! ����]�I"�0u����)��i�k���נj�������STi�{���ps�\]���׾������z.@��=,�"4��8@���Sh&m ���[4���� ��sXɳ[4�؍���!dT0���0�a0� �a7��4�H}����J�6�5F���g��$;�tuLUC�u�9�e� N��H��S4��:��(o0u���&��Do�1<_�Kg�cDm�w8�&�C7q���8v`��ɟR?ѽ{��̘L=,�����%?�󨹷+|F�޿��N`�bq�#��.�j�H)��-\�����Ĺ������͢� �� �1\�s[��j�;=����UW�X $��fTZ����s��+��G�0p���޾I7Zy:BI�	�aw�_#D�l��4yʿ�
M���-�k�L��}J��_��-�k�i�ڛwS�;|���}��RF���5�n��\) ����<����=��J��Z"�$#���YoV����G�H����99���h��3�ږ;�H ��Dy�����`u�� a�E- ����ģ<H�hN�`X&xϱ����?S���A�֩X��V��а� �E���wdN�.U�����Fpߦ�np��w���1����0���4�w�`�H��X�oa�I��;n�'U;@���#/���-ܮ��`lʙ���l�R��?z*�:�?h��Wu� �I��Ƈ�ћ�m���(9u��:��̍M���~'��� �!J��x(m,0v�^e,� _Bu�iǞ�
��4���SF��Wo3f�����N=��g{��Ba���`[x��D���*�ڹCfT��z���6���)�6 ~,�����.;%��Ln,b��ڜz���ILm:`��P��Vk#{�*�����6g�Qs�:p��B����7j<�v�e��ȅ�8��yDY��`M�4�J�0\�ͷ,��ܹX{|��������؝V�BΆMFiు��72V�N;%�i�!n@4��lε�>3U�+yXK����^E*��� V^�Kc?�(�cm�s^�1*g�0>�ϵ���Gc�]CދN�2Ƃ�uO%��
���Va�ߙUCޠ0Z;�����J�%�|Z��e���~�
K�����x[Â �^х������QmP���1Vd㳏+�ZuE՝3��2ˡ�u�w���~z�����Q��D�>���h+�}����Ǫ]<EB-�z��R������;v8	U� ��+��P�	���헺�:�J��ak��?�,B��6���z�6�-4:5���5el�j)��^M�5x�
%��N�ݤ쁭�A��õ��Vs,:��la7:�ι/���C��23	�5̖���ÿbK%�ғO�E;z*�	��IQ��@�"F&wPN���z�tl�UР�s�)v��d�L!���$�.�9a�h�dy��t����ʷ� s�>��M�*��VX�.ё�<�ñLO?1�i�hӮ�\8��f JUG3@���®p}����Tt�-.=N������PD	�4��t��R�b;�G�?��B�<���>�D��`�]����M�W+Q�f��qܑ���#z���N���\cjz����8����>�J3W1Odѻ�1{�ض&��Z�p��u�#��'�z�NE�!l3�¹>�k���.�a+m����b��Í����Y �V���4q�{��o�bv�W�!���`�x�co;����VHn�6��ٹ�/��,����q2D9��rί~������Ӑ�F, d��ٷ�kM�ܚؙ�^��̩���UR���\���%Jh]�;Y=�>t�$L^W��]�����}�C����-��Uc�F�����x��/�1�����L�-(��tsM�OZ�����Đ5�����؞��{,F	]�E8�0���s��z_�!;�C',@��Y�,���d��ɾ�N�S~�:���4���)$�� ��A��J���qYj� Q�g�mϩ���Ȁ[~���ͮW��o�ݩ�ڹ��2��uކ}��O������~. ���r���Uh��lgp�����|,���h��u�&(�_n+�4R�,c3���d��qAP�X�Q�X�(l]�`������.=�����e=�vʖ�e׫��k�Qf��iҷG�,�P;��\�?����%\�s��M�K�f�1gE�@��Yf�] VY7��ܫ�R�)X
mNV�T{QM�{�<b�/}AW�A�n�a��*�OBL>L�ĈY����R�hP�PKi�Pa��6��{j;�b�9�Y)�c=L;n���m~��i)�]~N��_>�֎�EG��ɠ��Y�E8�zLϔ�G��<sl�tݵ!
v"P��?|V�κX
�Xd�|�H>wGl�Q��,��!ڌ���]YHkt��
^�47�?�<�����rV���l`���[E�ch@v2F���mTM9@�8��<��Vb+��X��U��������|{�9��,��>F({U5Z��=�g������2;��1E����������n�r�Z�-9��z��j����=��`��'��֗�>��Y%x���&
�� FfemTa~zN��.�K
��Чs���p��of
�C�(̚�F�I�5��Vv�mrn���#df1�R6�aa|H|J���,�E���VH��'@�k���p�3�g%�͆FJ}0j��Ѫn�U���V��fj��([p�E���^).����1R%l�ڣ	��lj\��p���h�Gspe�t@�����,�P������z��5�3��ě_�b;�q��d�8�ml ��M3����`��uU���q��S&|u���0f_�M�|���Po%s�ʣ���a�d�c�yMF�`Jk)�v�����	�Sk�{��G1Rԛ*��x]8J(	��3$`�L�ڢ%�V39{v�l�}B��&�!*�W����߈�@���qW��xX��}3�eb�B�'q�c����yf�Ƴ��`Yc��A����T�h�֏F aIvar����S|E�8�$ՙ��!��M�b�Ǩ8�cs�02C݋`"oǞ3aY�L��j�A>�6���������z���Xte��jD��ldL����N�5U�kjX$�s�C��d�V�m��%c�#`�K�8a=P����k���{�k��q������[	��jx�C��P�5t�E�s��x�e��̙�a�SP��fk�kR�k��a������r	?����gzD1� ��:�we���lg��&l��� �ˌ�0d����__�xn@��-f����+-�1g��1k��qc��	��.����Ve'�0"=�|�]@�yX#���� p�W����*��ԅ_�D���±�G�a������/O��A�D)�(�Yc�� �)׸{�毰8j�N�\י�]hZЩh7�Q�$��1���î��qe�SB�~��=� B�
6K6�Ƿ@��oA�<)�R�.�3�g��:�f��V8��� ;P8^Kǉ�XF�ڍXZ���z0I�?�3����;�4w�UtP�`�5;M������7��/pk@��0PE�� ��[wӽ��0�Jc��!.���u�d��8CZ��sG�ٵ��%em��I=��%����I�Bjԁl^������)��w1����Ћ>f}j.-��np���$�=t,���7-�,���h;��ܫ2@^%��=�aw��r��''�X�vWc��1�lo����M�� �R�k��c��|�bH�ðpIPJ'T/zk���Vҹ�^O5�a7��J�k���8�U��v7?�uu�N:�ʸ��g��n���n̽���'+s���`�8����"^fQ_(b8Z �jz�:)�=i�b��J�ǐ���o�����'�E�$�1�	Bk�P�Q�� ��|.6.$�O���&Sf�Sx[�a�PˆZ���L�^�	����<NԆ�mZ7!�eW��=Dץ
��`|�g�t�t�[ڄU,�FC��D���^��5~�A�Ř����gɘ��:e����c��T�qL9ka�j՗�!�ռ�gDp��UKٶU�&L�F{�]��+x�l#&��B����+uƋD C�a�L�(������Ug��s$���ɱ��X�u;�r0=E��6A�+����<dO��Z�:lp^��/�i�S6�{l#��p)�5��.�?pԢ������8��~@F�9]��7)�b,�>m����,KoQ~��'m���Q�����0�{删��|����ν��1��<ѰS�{�s�1���c����h�丛��Ŝl�]U|�:r]jK0�sBE�\K�ly/�z���*��@Mv�q/��,i����v�t`9N%)�a>5�x�:瘃݅���R�%Ԛ���Ȫ��iP��jЈ�1uA9�ov(��ˏݛs�:���0�X���ut��<';�L[_��P��v��~�Q��ښ�BAv=����Z75��L@���G��]���"SE�S�Wq��e[A |�E]@�駟��C��9��'h}�_��.=P4c,��[��x��)���
����3���_�ɳ�����%��GK�,?�Ϣ�:2�!�v��'O��������=�qZ�u�D�R�����;�7�]Z��|B����xtn>�N�h��a-��B�C�n�4x�bB㴂3�&z'5L������c�[��� ��E�P�A'RIC+Jm���{i�RR3� Wi:�V(�TR����8�&�\{}g*���su��J��
�����	�m���+��9L�X��c�DE`H��waV	PѬ�`O�^҃���{`YDZ�v*���HoR���]Z���?��5�)�^K��"������	�d,�$n���(�u�=�ǜpG;�G��P8w"���&�*J~U�8߾�6%]�a_�o;S =,
��kX"��?���V�=@��>|�t�F(����t�n<�Un�T�`I�h�<5\a��kF`���_��v��%s�^'����4�U�}�~���)M�a'��z�Bj;:�n}~A�JĎ��\����óg����Z�a�kVOY��c�Y>�u���gܽ��W��1R��� 	&����Qr���DiOf�C�A�n���VC�	�Z�L��Q�k�NDK<\Kh�����9¦����G�-�>��"��즅�>E�9�9ӯ&f	�`���e��,�,Q�`�K_4�Gm����s��1����bK:l��d9%af��\��b~1W@#g�ʒ�n����v{��j�1hW�y���5=�,e�sǵ-��H�$@�s��r,")<�=�1����Ȣ5�L���&XC�oI-X�}��2J��e�*c3%3E�Dt�e�[�Vg��=V�I��Cx`�,ʌ|YY��Φc���O�#0P��򢝌�1>`���`+��Y;��ι�yp��� ��ڎU#�Ȓ>�/A������&h���3�NĠ���r��0�s�A��L> �Q"^�n{��o�3A���]���ȟ���E�1��1L�`��uҤ�}b
6pj^��c�@-;Q��૎	�(�v4�uճ"#�cn���A,��`������X���謡���r\�8����[�g�`H�E���R��O�`" �*&~u��8%������LO#�e��Ӓ��Җ�4���g��-x��+X �~3{@v����o-��V��i�n�������$����!��A2!����v�Q�J0>��S�r-kW�<s�4�:a
�>�[�jg`�������l����,pU�a1g�� ���T�?T���n��Z%��ٙ�-����w�<�N��%�:>�_�h���^�,��ŋ�w(�u���׈��m��4ͳ���L��E�3�Ko��ay,�l�_|1�����b,!L_�Q�GH\���m:�j��\�~`�����4��̢��h�;�Y4���zhu�`q��z��a�T��L���LV���Ј�`��X�}��iV��V�m���O�P;e��:z��kM3볩��'u}}�4�q.�#��T�8�My��~�݄E��u��[(ݤ$�Q;����K�W�����A��RJ�����o�*Pݤ�d|/�6ϑ.�e0��h�j�U�~��V���K�Z5�a3@����6m�w�E|��)c�!.�gi��a�	���Վ~X�>Yǭ��(m�p`+ʷ�P���3;
uK l9ˣE�1ƈ�R%c^s�c�㰻֓�v�Zh�_3�ש�k��V`rj��6c��M���a�9��n+���e E�k3�KA��w�О�%+ʎ�m�/O�+Z��1�Z�U�U���5�b,s���_����+���x���%�̼�h�&���xp��z�[��d����0�lr���f ~���v�_�p�Մ�nDdN�/Mo����K�ʁ-SF���L�WJf�s�Z.c�n�ѹj+�6�	Ƶ�]�VL-�)�q�Bn ��L��>�eu<O\S�?EƾݚyuA�L�Wf�l5wS�q9	� �PC�C���1�d��@py �(iq^hE5�-T�y��:�5�v�Y.`g1G!�S=f�/}AW�A슶�s�e����� 6{Ɖ堅0x��r�v�����e*�yG�¸�����A��c�b	�ݦ�z�sܙ�S�x�О���tY��ױ[�2�ҏ-��,8�`���dDX����� �l`��.[�Ox��U�"3��'h2�p��A*���tPv3�Ī�b�.�jI���DT�z;��ü4SF�~�� ĶP7�}�aZ�3�E�I���[a0��3�C�B�B�:X��ڄ�C��<����W(��!7֓���P8�s@��7�r>-�aFR��9�c&3:47v������;���ۑ �T�w��
)����9�o������`��������){J��Rt��j���X�� E�~�Ss� �V�GG%N���$ǣ_�<2G��-���� %�.75ף�q\�]6pi�yj���Co4L����F�y+���l�"z�E��"l 6����41F!"�٧s�Ac)r	&��ED��7K9]�S�����Z��i=s2���8��J�>J�h���Q�ʧAy=��1��.@����W'm�[,�j��H���
��+����W��Yz�	nW��Z�{h�EeUP��dO��8�Q�3�h��f����P�*eh-<<µ��W�<�w��}�1��Fz�������{���w������i:�G�<�A๏X_�?;�&�31>X�"���n�����[�mO"�nxʠ�4ΦJ�HN3.��m��ǟ?��!ĬĴ4�����U� n��t�N�%�чa�l,h�Z������y)��\�و�C�p|D�z#n`wH�� �����Y�K�x�Tb|���x]ˊX�����"�@o�Ҟ,V�����x�^Y=�c��ؐS���f��37[�?�cX������)�7c$;�ﻘ�,4��%A����(��?<ٔ�=�N 	u`zez@ ��5��4\��H��4�@[�-g��[X�$�aHl���l	�Vy~_�h�J֪��P]�s��o7X��nY�{h�HfY-�#��ݫ��/c����
w��ҼOt�<��fnm[�Yf�p�������G} F�Ndgx.4���K�^�{�B�"@9@�`]j�� �uՊ��r׊�ϒ�87 ��e�<A��e?�v�i���.3u��U-���5����<����ڀ �ۙ�-C��h˾�֐���̯�W�ew��,�G@����<55�IÆ�Y4����f�h�fj���dN�!r��x�'�Y���b��a�l7B�o��C�"M��&A �D>�%7���U��PQ# ��]s�V������<0������2YW}!}�x���yL�=A��v���i:�FIX�N��?VK��`��^����x�|zF�w��9J-�/(�����7�.���"I���Z�D��Ԃ��6��#C(�Q��F����F�OѫW ,ί�Ű�8@���	�����ܔ�lÔXN_H΍�,- �o�0q���E� ��' ��V��OiI>}��;q�њ�͢�+�K�x3nd�Q�cj�.��;�R3���,�����Zv��S�Ƅ?���EӐP�}��{�v�������Do�	R;��XZ`)�)7�i��x7v廔�^�
�z"=Z{��+w��̠���M|=�2�op�^0���E�9���������̷J�[��@�:�~�����)ZҍU8AKzѸ��jZ�W^���z�b�Y^�=&|�b���ߣ�v�,U��D��	q�\%%Fv�'ΝLJ��n�������{x]�w�Y�5���m�w.�0���$��Fcm1�aq�z��C:�n�k|s��OhN�q�^���J7��j�&���&��!� ������ҦLí��G3� �bg����u]�k��z9���(Y��\>��\��{_`%5�tqc��#���X�.�
`	p����RJ���қ���jS�wA��;�V�y�2Y��Y�0U-섍F�K��+e�L�Q2@Q��tCQ����e����4�s��:�LDj9����D��L�vV�
 �e�}��_0�>*<u�ٮSbp\Ɖذ�9����Q c��P6�R��}�gX .�R�9��>�JY�a`��	ԣ͇W1<�8�uҔ�k]4x�w������bZ2�4�qĆ�36�����2\H��F�3WW��!g�����˹XB3rD���pdRD�z��������?~l�~�tx���B�1g��z��<����E���_��1y�9�OԊ����]���jƠ�g���AE�+�E���=�5C��;�)D.2`݉X�wO�&5�sp�0p�hy5U d�ih�y_��R�a��bT��{=��N��,V*q|�'�XT��s���^c��ʔ���,\�`v��`bX�i��Ɲ���}BY��bRgt�'w�v�&Z�oN�L�N���x����E+�l�&�*�i��\AuC�.#�F�X���Ƒ��Q̮�Vt�#���oS���q��R� �&έ6��K����?�L���Q� �0��	tn=X$�� ��'ʊՀ�:X�:G��!�$���E�z���	LGq� ������z�U5��'sw����0l���.����
޳�E�?�ELV�͢�Q?���06�oܤ��߅�Xy�*��8�+V�� hhzl��GP~����ZRĢ���݃��g��8���&3A��9��������T��~)}�˟Q~�C�C�yN�<�b�YZ(*6�܉`z��x��M�n3z�)ʍ����`�K�N�f+�9�~t]��1�C,���Ă�{��KM/*zә�'��I�}��i�+ǳ>J9R�q��~7Ĳ�?�U��̬+c��Z\�	�9�t�5��?��Ё�����j'��Cvթۤ�H�U6� �m���jzP�^�޽�F��Z���Y@�=��y�hǦ�C\�.��ʃ����XL�(�ڍ�Q,- ��^���,cY����* ������i�����*)%���긐Ud�.���Yʪ Dv�lu6����y�Q?	F�ccB�s
zۨ����)����ᑥ�͏�?g�E��_�
Ť�E0$�%�PKQ�Ǳ
�ű��� R��07��5�Ӷo{,vY�o�2L.l�\�eK��S8-sv��3�i��Q�uN�j�:q��!���e�!+�{�
�[j���Es @�9S��/S����;��B<-��*&��/Z���0_TS�[f>>�y� ��xv�h��]�e����4�݃M��V�n�*~�V�F:8�Kf�q���Ǳ(^+;���}���:~{ޑ�(��oЈ�IM�끀J�#��$��P�<��3����ׂ��y���-�����'�6 P��A�͑�)Cޥ.�߂"��	D���-v6E�������w�:ك�5xP+�J�U�"0�Oz�����[���/�~�v�Snr�h��2z�ko]��JMנ���*k��zE����:���by�.����,:�0)�֒��]x�"��!];����Γ�$�� ������ʥ+t7-�/�ͯ�5M�YU�qW��8�U3��)S�ճ��b����D��[�&vԂ�2�%˫����4��c��S��K�W����*X����ν}9M�X���D9��Z'��}u8Gx�����>M"��iwk��&����O9<�b7�]?L`*l�
�<��3K��v����*&�z G�����������_:ڥF:>�aV�^�JVG��7�p,~,�t���; 3��D��z(�h��Ĭo�I�wzϜ�/�P�{��xH)��b۩�gP�����4u�n0_�č�8w�s��O[�����g���@���lM6vx� �����i�{����9���Y�U#�wm~9����<L���Ӕ�j �or�>,��h}��<S�e�9�i�ª��)��Ow�=����O; `�׸��ѷ����֧+�D�$�D0os��ICm��{q`81K�;�O=i���x��Xǆ1H�>-GJg:��Sl���-����� �j�V�>�b���'$St,�d�ױ�B�ɿ)��s�1h�c���f׎�U��G��T	��@gsE���|[:����� �Wޡ�9�矆�t!�7:q6�m��H����L�{S�zJK�gi���c
�ґ 3L�S�;��lT�IE�B�ol�,�Y;�j%�(��^���W87�����
͍M��8�؋�w
 ���e�v�Nᲁ�RZ!��8��.�lй���=ҡ]�&���^E,�Y��L��&��a�*��pV�p�o=N��%�(��!��ejF�H�Ch�".�Dv'�o/o>Z�S�d��"�j��n>�i[ S��7�.�*ގrX��dU���<{��'o�X�L�1ru��o�.�M5�X��V{	�u�56��N��A6u�hK�Y�?jv�y��M������z�&݁푾�s�]m��Y%��Q�vd��Xۮu�r� �F�.]F��Ho�rR�~;`ܡ5�pw���vW(-o��	eR�Y�}�������]��A�d7<��b��h���Z�z�
�MJ=�Cd�Kң�R�m�Ք�N4���b��o	�1G�LN~�v�F؁��	 �Fg�����_D�D+`n��b���:�l��dg��Ln�~.�Z�,�mP��$Y}�@�Y�#D�J��50p"^hN��)�Z�I���W��9��* ��O�|΂�D)�-�E�V������S�ϧ��x;��7~�'0&St(�h]���m�rM�n��y�n֖'`$��i�<��}���Ӄ���o�.��٧ƿ�y5ĉ���X,Ď|&��?|�ja)�����i�f�+וK���Z1H�
�!�_O?�����Z��y�Ԏ=���ԇ��"�t0�>�Ă�@ku���1 �I��1 .��v8�3G���S����6J�<K��d����$vBc�gtXpf�~3�N[�����on��` �~���)�-/��obL�!@]T�.:�f[�m3Ǫ�������Џ�����h�b� T��q�z�2�M/�*,�b}�@۸��.$��{`�V���Gk�!h�Vn� ��H���5 �M@�(�ϑ�"t�`A�Ek`��ᢇ0j��(��	K�ﻺ���F��h�m������Tm�xq݂]	��1�v�����u����*qO��tz�6�%��.4-{k���,�2��,m�ƿ��MYb����rtA�?돥'���圫�Ia뾿#��=ڒ:1oO��;� �Ђ������;͓�]��,��~�<$v��K���֗J�3���c[ [7~g����h��w`錭���c�U�+N��c�QD $H���g��e�v_q�}��I@W�k�J^c9)��� �Σ��[X�l�A�U��&V������l��f ��a��[����˸�; u<o����3Ph0��}������s8Ϗ8X�)�u�Z�%����O#�mt��(PE�������^D)�����S��*�N-�zN1��@�c�pb�s���o���SN'��H&��'��	���X��L[��Ev�˰+��ۗ�6|z���N���]}J/#��/l~YJs�VFVQ-6���YTu�5Eٺ�=�	�G��9������(L����5Ö���&r�\T�YxX��P����g'M��p��vJge��g]�~�A�FS�b=z�s���`�ͳK_�4����E��Ejy�����'���*�y&��g_�=��<��瑚���� 4� �Zb5��]vxo�s._����,����Q8#$���3�U���q���>%�u,�)J.�a)
\�ZĸݧiP���R�;�n�ʾ��o��`ilu<Gt��\����ӧ. ��	��ܥ4��GP�k�X_$��\N�Np_ۑ�M��$�"kK~; �	ӎ�<lA�� X�7���+�sZ�D4L�Pgꮾ�����}�x�B��Fk�k����� �۔��`7(]���I2>��[7�k e�yo��Զ"2��!� |-C�Sýk��������O�1\�C��{/��j���j4�<([Y���q=����GǗ �m��&ό�۞����X�8w7 �Iww�~�Rz#���חmS~DO��·������� ��F�o�v��*��lFV�}�v'�D����/)����C��N�s�6~�I@]�O��ln%�Y(�V��Q[��gy�o�1鵕%���Жfg�}���\�⠧1�/ۦ��6l��,�x.�{h���)A������x[.�0��p�D���13���J���2VVj
%R�Y�Ա0s�p)k�� G~l�d,�9�m ʷLT�|݌9�eGl�d�db"G4�:&;Kcq��֍�!�>�[�?���d}dҪ�p��%1��]�\W7��������� ���J��]l4?�˷ .��X��|Y�Qcd9�X�%���*'g��N��j�!6Nj��tk�趤ɜ��l�yk�{���bg�q>�\S��2J�t�i}`lF�P�\/�1$�pT_gH����' tCi�n��pʍ҈�^V�3�1�=4%���wKd�+x�>���v^ĄWȀ��v\�ά���di��X&�V���B�¢��@Y��Z�N�O�2�mv;L���3�j؍F�$�i��S�̌"�U��t'�	[QA%�j;@a�{}3�ő���D��v�@�|$b׵H�>�������F����?���q��>��
'� �;L��0P�����g#]z��2{��-�9�*:�v��5�#���P��"w�O��}:1K|��d�u�s�֝۱{�+��kbf���W°P�����__�N�u�i;�n��m��yCzr�k�3���N����:;�6����E�Ul����K�`	d�F?���1O�Z������K�$	\Ew��Fz��<-�_�����Ą����1O{�$��s��K� ()�Ow�x��>�l��EU1���(;��2@ю�}�Q�a��U���+�m��I�����"�Ft�!e3m�CD8�V�P������6o��\ͳw���������s��T=	�X/�ߜI�Ϧ�KE'�F2��|�b�9�x ��8���wp��F P�c�cV�_M)����U��a�����SJ�K�/0H�N/�>H�>M���`|v8�	��>�{�8>KLL�˗3���z&.XN�-L��g�jJxo}��`��^ރ5��,t�۩t����"�����"%~	넾Ԏ�Y��`|��G<+/���Ʊ^EKe��!�o���7�fyo�:J�2=�:1�^��.�Tw�,F#h��">���"���0&.� @�,�e�d�:���1n{8 f�g���ZO�����	*�;Q���amF#��3,��4QPTb��ui�;��w�B���vy�]Y���?۬��"�!c�r���o�=�se�7��H݊yU��s���S�㽓�Q���j/�G
�c�O��󳃣jd���>�GkFG(�$�(La�a������!���������|Y9Y���������k7Wp�V@�G+W+,|��3��.v�zmuw��n�M�����ƕ0�4�ʥ��5�Gs�髱B��hK�)|��] M���"xU{�Cp,#&@�I�~y����i�˷쏠�
D�K���l�f+x�Г���`�zm@��w���Ĳ�&�{X���/����)t<l�����H_kx��@�7;@5?,�N>̾�6oW� E?B�*:<LYf0T�m'��W'�v�t1�Y+�f����dp;Qȱ*B���dw��&�{t̨Sx�ߟ�yeG6Ė}Y.��rx�]�����Tb\�cT�`�D;�%~6���Ʈ.�[jqL��x�(a4S:��c����-�1U��I����γ{�x�y��_Ά)d%�>o_�	 ���q;F?�6ô�y��M��-�d��I�"�#9x�a��wZ�9؉."-�hc}��@�x&��}��uJ/�h���W�:�+ua������]٦#M�� @��f�VX���3>�A�ܦ����T@�T{1�����ƗR�'�T����qA�h+�:2</0}0 ��>���i�� ��6B�{e[�!����������4'��͉Y��6�i۹w�2Q�ukR����]9;��1Wh��ͽj�{X�}B�yB�>:�*�K��dwKy��QV�v�mΝĨ����W��������}nl�kL��]q\�(�rܝ�5�/���<<���v�݈�k��ۃĔ��W;Ƃiy|Kgj���m��;�~���^��p���rz��-����TUn[i��&=W��,ژyz,��jn��
�3SQ2�9����"�>_r΂3�,P���n�[���qZ�:��e�X�c�K�E�F˴zme1���.Ȍ�tqN6�*�"Yݧ �*[��6,�eƉѰ�b,�c�;���ZhSJ�U��p:s��+��X&����G%�G�#u26%D��>v����\�:Wk波�޻�9�k���rx�P���ω��s�_���s<;�� ��|Ҧե�4�.9�3/k������	l��o��q���%�o!Ni&�:4��l̜��y����� ^�JH���7uO��]F�9���nk�!`�pb�6��Rb X��g���i�g�j��Ol|`��<%q�$������)�x.���T^q牢�!bWK$ ������̅[������K��������xm@4p-\E�E8F.�l��V�L ��GI��ΨʹƎ��b9��"����4�b`�2��*ie� E[��8����m�@oF3"�\��B�΀7��ܭ̑�Y(3N�	Ѭ%����m�NϦ?����c�	\�;���7���������O>�\%_���5!T݄Q�������T�/�SX5�q>?�]I�d�=��v�w�;�͸�~"C'����qZ���s�������o�x���#��`D��E)̭�Wt���#�}�����	�Ra�&c��N�?�7W����h���V7-�t<}���i~T-I}�Z�D`�H��&��؟a\�;�<k qYp.�55;ڝ��%�tʹ6+t���6\d��]�7�#� ��(�lB��ߺJ �����H�g�d�IS���ѯ��!�B�pvC�~s�,�TQ�3Z���_�p�����nO��Q[���wߤW�n�ޘ���	���G��&e���44�����In'���e�R�[L�k3 s�{�Hn����� �,�V���H��7���х�?! ���\_+`N8��`��1��~=]��_� |v~:�>Ld�T�ݫ���Wig����q/�7�ΡZG�ЭK� �V�iʋ� c���9�>
Ķp,�Z�;}=ur﫰W8�f��ҹ��{�[w�C@�e�k$���A��%�1�3��D?�G��qV�OQu^D ��cvo��p#$+[ϵ2�Uۄ�	�}m���q�D�k���
�7xɬ��r�	
xa�,��� �e|����	�eNV���iv�N4�}��x1�j (!�����!�f%��ļ�+b~��pTvSĿ	���4��)>>?�0��IC�Z� S��b�KǲSڽ�W|��c�ɞg$^(��)���pTZ���4;��l`~�=2�ZCBٓp��U��(��
��\[��-���< �R��|�:�7ëD�aK�<7��漙^����zT����A��=m���N�����^��;rp�i|Zw{S �r�2׷�(�
_���un�q誅��{��ahl�f��(��16�k�� ��>D�?�6�
�H�E���N>�E:fs�Z�
���d�h����r`oI������{��x-@]Re�[�aڣ�.�;�X[vWĀ���3�Q7d�3���/��}�3xXԔ���ie�`+��a�s�F}��`u�X0f��f�+��R3�@K�9�ߛ�0$�6m=,�1cD�A��.��Fgf���9�-#�}NL�$T�_]�&�7��>���&F²�����,�л ��J;ca/dKF>�M�f:I.T+J#-����B�C�ik"_�i������
!��7X`�q�~;�|��*�۱�E� Y�!4}W���"�aA�]���hܽ�yL�κ#0o�:��.�<��߾	׵|��r~6����Jx�,~]�,F>�pG[�s\�a��^�,ڕ=��O>�l�p�ס�ћ��V�YL�ȳjl��Z�U���P�s���hyN� �r�Ɗ�\;3��v�0U�/)��~�Ī�n-�-�6L�nP��F�H� M�Z�M�� �0j���9Z�m�}6�V`}�֖Y��,6 #�}ų��_fao�)�+�2�׻P8�Z���'+�	m�,]g9�a������d0I/�2�8�`��ϥ�����;�>�mph��/p��ݹП�BTH[��hʵ��?���g�H��K�V+[��{K�ߓ2���܇���'�а�S�|��lz���N��S�"�6�i뛔#�ǉkA�_Fpl-�9�kDl� ��#�G��u ٪��l�az�h���7��s�q4�D�#k�0�q_e9��"s����,��Q���I�&���V�(51u��r�M�)�z))���s��b)n����$�g�@O��:,�!1��R3�/���ѽf��f�0SXʊ�IF��"nɅZU��=����s��V�>�b���K��]��c���F��Y�� BR\݊�������UZϩ����n����U;:��%������ғ �4z�u���\�ހ E�(���r��X���M�g�� �Ӑ����Xl��<��#t ��
�}�5������<��i�򽦍��o5|T��[�̃l��{s�:�?��"�s�y�4�s[���*��-�	fd�C)���+X��2�G�bI��"�v���L�!g��:Ne�����WPՅ(�X���� A�O�:�w�6�8d�ٗ��R�~���J4������+�X��H���1Q���3�	a���1cqJ�l1H��g�n*���� +Q��0����h�V�M���I�2� ���l'<�-	8Q���g��h���g �߰(��[�[�I����t��s�j�������g��t�̠g�__�D���F�e'ى;�M� (�<u�_'*���v��r���PN+�Zz�B�#���:�t�]p�0����?�yZ���v}�^U�|�Y����͇iu�ij8A.^5צ��r �������a��n�%<&�X ܁�y�q�j�w�������L4���q�m�������ۿ�y���T����z&�:���)�h%�=���L�^C���qӶsj��l����u�t�ϒ]��(۝>PYL7��.U�|v�a�������%bW� �D(-�`g�����á�:��w"����G�`B�I��o�S�2��F����(M���Pu�����+�Z�����N�d{i#�^��~�/�E�0� ���&�Z�O'��	���ճ4��A�:#�Q;�_�͗.�WOp���oig�E�Ciw{����$�8{��p ��c�%]E7����ᯖ)ԡ�P6r��tr�s��o�oa��ya�x��]��2��KʄO�oq��t�eA:MH�m﫰��K��)ҽ�k�67̸bѱ�r�������&-E�S��D�cw_Β��(v�6�¼�2���r���%q���7��CH�t������afy0��d`E�vl�|���g��������5s�>��01�d�ce���+Z+\������ЎE �Ƈ�Ǉ3>ǧ��s��S�%n
��cN��9����j7{A֥�TNB�Nʲه�\��%��q�k�k�th��rS�{ʼ�>y�7l����4Q&�dڈUH����B�,϶��˔l1U�Z���>� \�����E��ky>�ۍ�i
�u�Z���7����p�2Q��3�3 �@�������0�l����A]1�ݻf�������X�t��:�����p`7�f�����k�s������l�h���C���_?�x-@PL0eek�9z�e��1�j�������Q6�A�uxQ��f]]G �v^z��������wӝ��2�3A��`Eѳ�k�j�`p7 -^'�`��&�8�D	�؁�M:�L���NX�c��ol� K�fԷi^b�<F��+��|y���B�4�X��ff�\�3&�\)r�\�ӊ=�ve�!�~x��k�r�c3,��!61 �!U-A?姖7CT�8p��3g�j]�f����)X%��^]7��\�5�M�mN��'t��<�����U T�l������9O6=��d�.�,5ZM����Q�Ӝ����S�^��'�n�J���"��vx;�G+���5L�ң�\a��κ`�.(x��N(A� �v�qJK�H�Ͳ�?u�l�x���P�3"� i<�b�y ��r��@�yu5�'?OkSv��W��{�QJ�6ʁ6�^��N�"Ks{_���S�ee�K��!�I]�'�n!�,r��(A�Q�u�`љ��#�_�i� CS�}�99�jۉ����k����9���o�S�V;�52Ԛx6Z��<�އ���"d�� s��%��2���j�m��A��2;l���� �5�Yj*�C����v�3��c�������$�������)�M��~N��Q�LH/�Zpj��"eD�B7z����@'8V�� �_�zh�(�U(@q�I�R�%1;�"��]���2��c���P[�hq2��p��+�7lu0J�	6�2L��--Yz� 0�k��{-D�j�J�&�)�z�7,�.��(�̈]�����ew����1:�(8��ľK�{�dV� �WY�A)�R��d�r��ag_-s� ��?����,�+3gw���
�\cg~�Fy8�T2�XbSg'�&^��G�Fg	���G��~_�[Q�� Ӂ�C?��rC��ҮQ���� ez�ٙ�_h�b~����er���I��� 𭹪����1:	V�	��^�F��J�O�����R�rA�L`ǘ�<d�� ������p�e��@�IV���\���1 �uj'�-��\���C��>w�f�,d�^�I,�eR��&�@~�k�h]-���g���gh�	�!�p�m@����>Ա;A�X��z�`Z���\Ie,J���a�W���,vjvp@�2��a���f��B��Ţa�l���C��p !�S4���vU�d���3�oue"�u&:�^:y)r��#�r:�a�%�mv6��-�|x��c�������ī�dj�e��.���5=�X�@�����#��cȤ�Gҳ;��$;z]� }���hV�c���O���d�����Y��ЎG9D��m��P�?Ĉq#��j����m�Z���|5� ���˜��OG����К�&��Ə�-o�G��ui�yz�����R��a )yR�W��ѶX�{����`,q�Ͼ��ޫ�F�wX]�(u�]���; b/8�G�[4����&�2b��&���k�!E�\uW.BӜo��`:�N���d$d׋�5[��[�	?]I�0b��^�\7�&bW�6��������O>A���so'4X,��)*	��:{2l��B��J���-��s.�z��s��s-�E��,hYG4�@Ъ[�s�/G��2ǐ�Y���7�9����o�Զxn+D¦+��N<�.0�fJ|��\H����D���XF�����ŦW,F��þ��Ln��Q��"j�L��.~��Œj��s�����|����[o�{��X�>���$�������_���$�Yp �A��9�\{�LB_DK�cǗǩ^OSE7��r��h�t�{j�:a��Ӗ���Q��g�@)U���eǌ��]O�u�% Z�i&���)��8�d���	5VQW�����?�,�����b�v�?@����d�hhq,��R�"�+���yD]��ɶ'E�YG���U�Qۖ_�����c_�:r�Y�������WTY$�!�z��p�l
�9~|�7���.�VKZ�jI��﫭�*��hyD�������;���l�'�3Z(w��u�n.s��=�iG�Ӫ!"����_��>��7���ε��lڰ��9��X=s���-����v2'W6�'m�X ��W��rW���u�׏|�m��t����Q���0;>Ou�����2O��z
d���UEGYv��԰٦F6��uI�q�[ H֗Y���Y�@��_����bWU����6T�:�:nP� �a��wf��T��c��X&�Э�����_7�2л��<�hMͅ[����>��ý��O/����|�z&�g��R�Y��kO�U:�݇/X�|d	l���v5�~@����V�=~w+|�����Ĺ�;w.f�;_}����b1���M��+�צ��P�m�z���(v�uG�(�H������qV@��*�o���pƦ�d�SA�kh���}>��;�uؘ�4-��x���R�*&,���)���ҩ�l�B��/�,T��ݿB�X����i�!f�,r&���r���/��=؝�	e�9�i
�:솿{
=����<H˵G���[|1�{�K�h�a�g�Pp�r�eX�&�E:��y�h?�y7���i�z�ч��h�7�b���.��u3� �o�3�UFILÜ��Ll��s��?���=8_�{6i^j��l}�������!���\�p9�Ql>H�
a�hI����>(Ҟy��4 �c�bg��l;=$�l�.]t�l�Д��ٕ0�3�6���X@�W؇);u�g�����Vߤ���#W����N�1 ��A���&t0fP�6��1=��������1�t���=�����<� &Ac��7ks�dh�Q�[�<�}� hWPA�c.��w�����l�8P��3�v�ݸ�P�	�
B\�T�:�S�+�� �0+}�w4�"��w�������dOe"�O�T.���8�{�u�b.�щ$w�!b�EE16QU	P#��:�d��PU�ܜO�G`:*逬��C���NK<�ː��w�_ܸЋQ+2Pᘬv����1�ػtN�� ���q��\j��Gh��4*xV,g� 
-�
� %=SE�{~Gnb�l��	>��Rp��y��h���`��P�P��ln#~V�lf���j6`˔��a�G�z(064v`�(.����l����g�f�ݵO�V%�_�g��0�1mmk� S���EZd�1�����Z� ��Mʁ�&��3��Ch ���ƥZ�;`���j�"s,����{�����1<�G��l��9�H5gm�N"2.R��h�4 Ң,BE�J'��uw[)}M60�:8da�Y���-�;�.t�&g�H�_)�Fe����bRu��׼���a�諓M�fR�Ԑ�
;�5d�l/�?[}��y�#�q���z���"�����v�j0��L�W+
ֱ��_C�'���0^O���DO87�e����Q/��?�z���`��^���:��2���+���@�dtL6#i���&�-�8���};�L+��������EF����w�ɟ	����o��k�����R3�]5Mm�o�s�b�%�_�P�	LU-Z�v��4V<\1�5]�QQp]d!��q0몑�NX���^:LN�\£��~P��a���܀��� V��e�|���m�v�g`2�g���.̱������Y��ħ0k� Ν�rS�{�a��{��8��ɿ��QNx��@�R,]>,�Ct��{�����C�[q�F��4�68��N��{/��1�@|�\+؉��.ɀu���O5��zdu����2�:�ѽ[7�c�^�U�ۖ��:J/>���DyKI�X��@:������Ѝ	+Z�[Ġ�q���9@�\`�p�� uǱA��<�Z/��<mP9J1�>o���5�
b��J@7�Y?��>�Aw��	+
;��c+(V�������A6��X�m�y�� Pe/ k�������0�s�d�1GEvC�����OǌS�u�<ob�}V�ʚ/��J������+��)�D�`0nxa�QҌ	$4܋_��!k��oP�?��*���,�:��0JO�P���5��q�!�������b~. �c�{�����D�˯h��<CU�.�R]l mD��Q~�����\���8PM�25C�Y0V�8n����c����F�����g���DmW���&e�2@����:�W�k�h4^�ͳ��Q����3(am �Q�b����ŵ)"���Av{S�A3��󴊍�%>u� ���W�`Q���XEP�,���!��KeN~�yW�8>+�i��1V��g���~�+�:��-&�
�J�~���GP�����x(03�S��lV���dYa��#PqB'���K����.�9��v��P�˂�h��ш�IT �p�>��ݴ�22'f�Q��,~�~���y'&�G �i�Ma�>��8�X�T���oÎv@vRY��A�1��fh0:{ʙ(~�u�bM�C�bcj��ֲ�$���H��z����X$kة꠬�Q!�?�D􂈄5���<CC��P9G���3= )��ap)7�T2A�D��g�~�r�R��Y��@�~�8�}C�8wE7WTzש�k�Q���V��u��d~�8?�Y5LK+n�:d�Ej`W��΅T�џ�(�mC�O �N"�.��Z�����RWv��&����8�hr�Ԁ���@\�=�޾H��nj�3i��[�����Z0S�q����,���8�'@tx��%�,��+o�����d�u�脻��t���4�׳��|]�]ʱ��y)��_�1k���� �dK;s���y	���28�C����X�	��%�}��L���a�h�jз���4��~�Z,�6���`�
��W�#ّ	�<�&�$e�z�0�*	�e�u��=@t��A�Gq���Ct�����6���2- �~��kxfW �� �2TM�¢!{�_�� ���W��󚀆�Jgh=��)���"���20~�z�+i6|����P!gP����%˴��c���Y8�JǮ���~&�d�s
��@/�"��Y�V�G>~�`��sP�J�ӄ�e��=���ł� ���+��g{, 
�tGGl��s�@���0]
�t���ѵk8��o+;��Ǟh:Q;W���C��e� V�=�+���<�GT����]F+����ԹN�}F������q�`���5C��Vy�g]�-���ʱ R�v�$����[c�*�A�v�M��?�9 ���d�4;�n?�V Q��m^Jqٙ�r2���C6so�3F�q��������OfK�N���_����a����T��y�A�~?~�@W�A<hT.���G�s�uf;���:��VȨ9Ic�����%�]�#�ʎ�<��N �:�����r�@7�̾_��������Zf�J(W�R{��1�3B$g���D�0�.6w�ڹO�Y�}R��gjg��o�	���u]���[�L2O��X�^ag��0~55�����
�s�ea�fI�����Ca@�՟��S� ]>�iǿ@�
�h;���4Q���,S���  ��'�Mϥy:�� X��9�yk�
�X���'�v�e���i�/��T����ܴ�}�{&��4�|�qݧT'[uĎ����2#v��� �����B<M'�;�v��p��� \\�,���Ք\�#��� ��M�ݴ:��+?�����M,��r�=���%	�����l�_�Ua����#���G�ÿ�8Hc\�]���r���al���?|�^ ��^F�����t=ѪeG���a�c4e"?�}�3&�Y����0{�n��~?��m�a�v�e�\G<_��ݾ���Jw�ъb;�k�� uf�XWyf�(\��Oa�h�7G��	J*��4��K<���F��U���hDN��zN{��C�_.��B���(�La��
�iG �"��C��4\E�'� �kaҽT��I�\"ٍ����~���O>JOa�y���6x��h�153�Bς�u;�t>v�w�����L���c�.�Y@����m��	���&���{ϖ�`l��˱�FJ�6��y_;�v�/�:1�<�������Z�l����P@��#Y�W��c#&I$�ˎcOmJ��.� _�kf�j���8ۍ6���v�n,��\�jϹN�D�W>�[0�W5e�<ρ��ϋ����ĎUy�M�ctws5�Zv6)Q���y.4vLEɑ��!"&���.{��%�s*�í>�cz���@�$��<̋]jܓr����1g��%���I�ڳY��r:Q��m��&S ") �e^��R�g�>�j��,�"Ǡ�v-Z=t�ֳ�ک�\_�K�,��aPфn�� ��r�L��@�o,�'�o��A�k{+÷NV�燹���L�k�.�@8���ǼV�x��wU�"��p����
�K�.�Z� �ݽ��.���D �l���L��U�J�ْF��6ed.��-���|�إ�Eb���:�� P���=��?A}g��1R��Pب3�%*u(3�b��8m�Khuiu���������HvI�g����ѕ��vi����w�{~��;,]����gJ�Fb_`bB41s`3��{Z�w5�Ӄ0.�1M����Y+�qb�x9��l��1&��3�R�G�1��j`2|띴E�}�P��s���C�nބ)�J�sSi��y��4�j��A\۔����8W��dfղ��`�?\�0`�6HP���
���o�l��#�ח39Op�|�&e�m��^��6�������瀑2&�1��`��j�|�4��b�i%-m[ʫ��罏>����B�c�����X�Dܛc�?B��g��e��YK �
H蔪Dx��.[�Nݫs])ͭͥ\SE:Q2���t�k��?�=H5k ڹ6cic��:V��i����������[�!�@��cmw�����G=@���/�R�پ��G�,�CM,|��S�Ԗa���ܭP���; ؔ��,o�⎆	�>�q�Y8�X�^<{�F7%X,���z��n��A�i�b����76��e,�>�>M��:�|
�,�%�b�PP�ykJ�)�G�$��F��k� TE��ۖ��0y���bܡäp�D���?s\��.�v�9��k�D�TH�{] �(u1��v����c(�}|���MP����D��!_*��w���F���;����yE�{�9!�2XU?;�I#X�q���%�fC�K�ڙ=47h�d�����(��>ϲ׿\ (*�(��Qu�1Q��#��s��ʖE�&�����r��x��òe;ʖt��$l ��H�yH����1�-mQҗ��i[@3��9� :�G���>F*��]w��`�=V�)��aA-c�2�.��5�Q��ڱ�3���e�6[��dؒ�@SH��ef����?�6} U��{����on6��c����^� �I�M�9h1��Bǀ���c��v\D�0M��	V8��[��7�����M�Fh=�e2i2��A]`W�o�;G �iv!��5�)���2[�N���% ��`\��ĉ#A&�P%ٝ�b`:�m��&�d�!	Z'�=�A���G���2��^�Fg�]2�P�de �M�cT���ALN{H̦��&Ż �!��U�bz�� ����_Rz
�2CAq0�^�����u��� m����k��{��M]�g�]J5�Pz��y��;��B��!^ŷ7���G[�6%��#im�>9a=i���Q�Lg(]�52�ƛi]O��F�o���TR�����HZ`���[7�s/��S�Q�v�j�;0&]�\O�>�(��-�L�'�j*���~�������	,}2�V	d�w�ܫ �����5�uB�����1�r='a&�<�s�����X���-��Kv�|Uҩ���+�V4aP�Mk���w����+���O��N�1nl|��SfĠ��]:���1o"���)�bq[�i���Udq}u��&�f�k�"P�J`��Ug7%Qr��`�~��4e����*�ts�\��?�2-�I6�2%�i�j#��+Yk`��S˩~� �d�rl��_�I֚:��t\M9�'7��O��t�gY ������+��v��]U�;i��bU=�C ��TȞ{���X�=yH�
�8d7t�!�l����:Joo�<ܻw/}��OC��F7�"�JV_K��
`!�*�Z��� ��~�R������Wd��.�Uv	1�*r\2�����gT����0:2�*mm<k�l���κ��eKwY��!�I೔�Z���z �J��f�2�T�Z��s���Q���FT���fu���  ��ƱY���sZ0�g�����O��P�R��q���j4�FW4d�Ds�7Pp�2䶝g�_��ؕ��s�	G���l5jeX�7�pf�zV��0m��!�]�WI�����p�
ϩ��|*�Q�hƽZ%�k���4��X��{=[(i�\��#߻k�d+�1���IZ����8��:�Z����7sj,�1Ti3���!�je�*�5���Gp�x1tf���b�`�!�4��)#�C&�pլ�]@�Z h���(8�~7��<ʳ�G�9{t�r$ѦS�c��ae�.]'?~�`W�A��Hj���v=ٗ�s�j
qN�R��H�<��!�lqB�C�g%�+,��L^:;#�����Z����;��=[���1ޢ���N�Y8#I��"k�D�.�f����y�v�8��I�爿�C��v�!��PQ���-���|Q�u��R~p�xT7c�	�%��e��V��ɰ�`G�Y�B3���%4F� �Y ^��8��4T4ٽ=�����qk%�r��/�����f��rLZE^�|]�����vtlyL
w��B�L�z|�VM��%�*Jm8���R"�}&�ޮ��7X8�#�t����*�I�̫�oĽ����hT)�."l���䵋�zS��{�ΠgB�����8S��k3��d�t�]������>�Kd"���������[��,�˙F�]�N����0$�t�M¢}}���Bo�.���O��z�Pw׹��( �.����"L�6숻~K�͔��x6w���k8��g�T�������9@g�	!��>�=�Ce�F�範������J��s{�g?#�6��3�k��3���OR�d�E�o���M�z`w��aW`0i�S7z1ˋ
Wsl"��K���ڊ�B�n��ص1��r�����s��!�12��ez�����<� ��e�磔�Z㿊.@�ѧ�[º�W 혳=�X�:�I}��N�j���Au����>>��z��d6����5P���$c��1���c,��O�FV����U�_;��x^�-�]̳�S�Ja���|v?-�k���qԻ h ��Zݢ"�26J\"�-�|f4C��7��l�,�w�ˉ�>w���\�'�c>����t��v�Y�4v�/$�j�]}3G$@�k \�=+ӑ��WXm�-�)�'� vRi����� O�F���A;�q����Fx�ɴS6�]�V��UD���@��5��k��j�a`���q���ƿ\͜���G���Mvu��+�� g<!`W0-���3� >��>�)&�A-�'����pUN��n0�'/N<3�_9�5��u��z��X�z���訚������Fz� ��z��t���/'��"%���q��Wu���*��Mu���j�����,��"���1��fðCd�.���U��Sg2��k��ڀ M0��,��g�N����&����:Nq.���(oH�:X}�4W�F�ea�c'����߅��99���ўA�x~nW�t�
��Z��j��8��.q�����C�}����łW�����s�	��:��ȿ����9�f��?���Z�th4�gx~'aoܕ�����!Kr�9������5<,�q^�U�F�\M錅�mG#:�����F'c�u�_ǂ�A��C#GQ�����\���;�Laox�u"�i�P��Qs��b�_�Ԏf;���R+ i�?�F�"�k�{���0�%���^<�*�¢�>yD	7e�s�捰�ge%��$e9� �N��AG3�X�	���y���c�%���HMc��ck��   IDAT*u�i�߄��,h&ķ��@wT(��~,���� f	�m�N�-ZpWaJF�{�����g��q(}���G� ��=�j(QZ�9w��24]c�f�_N�mD�e,�3x(�s�?��>�h��`�JyU]�O���u�[\U<�Ӌ�����2��m��S�d�p��Q�pޕ[�M#�\C���gOϦ! �l�3��݃��}����ht*��x'�(�؍l�C��&�8co �� �=$�[���/�:-0Vl//'��Ak��7*`vt��'-y`��LYk��E�N4ݿ���e�2����?�$���|`3t�|z����U{�n}���L��|�eʇ
ʝ�;�vq���A�C���B)KR�ό%�V�� ǅ�� ������KbV��R	?3K�Pm��Ќ�:��*��W��#[kڼ�q�`s=ky��������'�"�b�g<��J���z��F�	�.��Xggj�B�(��B��m���V���㪌�1�ۖ�e����MѮͿU�{�

�^�Zxl�6��l�O����n����Y�%�e)���0'4�v��j7X�Zǵu���8���B� �M
/$��sg��%����4N^�|���yNys�c�7R��uV��c�#e];7 ��:(ޞ�`&���M�g|�YrE0Æ�0tN��� �k&����<w��p�h�(���g����AE��Dl�]O�e���s�S�T��t�������{[ۛĥ>�w]���!��xr�@��S�ц�,��e�ʷ:�����ƛ�Y�}9�2�SY���ü��_��<�����nuu�W��zw�u�C��3�!�����. 6r�����j��	�g)D���株�uwոL��4Y%�2avVo�:�����k9q�Spq��D���n�Ab���=SϛњD7����[�#3S��3���9���XW2.t�������:�F����<t�)�DQ8�x���N�v��T�IcA����)%��¢9�c�����=bk{3��D��ބ���OO��:�m_� ��F��#��M���(m!^��1<}�|���� ��c�X��l�N��;ɮ*�mKg����,��>��BB�g(�!��y�,4P5t��R6�Gפ�I�h-&���^I�燂��<į��Ż5_�F�R�S�R#Ue�ln4�7�O�x�G�,I眗��stX��Dd�z�J����VC�o�
ӣI�L�"��)�j�:�j��	�;x�)�'҉S耺�H��q%��F})�M�y:� l��`G9Z @��'�h��ϻ#�j��m������ �m��1n�r���O�E��x��@���6�w��&ҋ����f����3�S7f��<�C} A��J4�t} �n��H� ��hv1��km��������ѣd!�h��3��`{��q�k�Mt��\�y7@8n�D�X�Mt{Up��2`��}�b5��Ĵ ;���a�|�J�q�N��_�M�le��Y���\Z.Y�e@l=�S.2
���ώUt�x.�=�by��*���(�qpqqD�<�~<��ql���em�7��qRBU�b���C�(�\��\e��_�����y�'�����7�@y�`�d�dUd���4rT�".�A�YѵX�5�(Xy/�AȔ8'm�23��2[.켷�!K�u�q�a��u���
`Pҝ�kT8�e{}���x��}����Pc&p����f9,��]0��i��Rw5�c�^A�	���n
m$�D�x=��m�^@"x`W��E��El8A�Y�%�u��r��~]�ὤ(����b�pЖ���ű�^$͞ X��M���(Xb>w�;��^c��gK��\��fɻ�5��k	Ǟ��3q<��[�+Ք��)k�)��Ї��������ҟ]��(gq*ٷ_%v�`C��N޻L~�k��y��չæچŚ��W�}��|�}Zt���zm@�=G2)�$��ENe<�!�c��oD������}�>6̯ڈ�5+�+�xP�k#�r��AwAjh���������3Hy�,S�.&sb�#\T:}������=�>��z}[t�6 ��X
ϣq���o���ƶ�o)�8�9�#���W���B}�ʎY�9J'�,�u|�ۈwW��L�ؘ��{�|�h:��aw�v�f�{X�-v�˔�ul�#j=�-����)9	:|jtN���W߼��F=t� �ݘ�X�lPf�ڵ�8���Pm�	��R5�����)�I �*��d�iXy����zz>2��1�����ӧS�� �s9������E�cr�j�G��`V�[�<�:�3�ҩ�ci�{��������B��7�a�Uj�ѯP�2 ��������H z���,�<\��g�C�v�!L�x]#��>���O�����K��� �%���7:_�p	 ��~3f�c�@��l�9Ǳ��kG��1w�hL�xNN^�$��Co.�����+Ԝ1�iԨ�t��$_[d+b`X���y���M/�V_����M8	x��.���딵�i�q��`���q�ԝ\Ǎ[�O��9_��`1�~�ZzI����'O��2�tnr,K��g_��J�hC;;x�����,������g�a�&��x>|ea�ϥ��Q���ؐD�C=�����5I�	�լP�6Z�3�#
�̻�� �����c)[�(�p�K�r���a�H��a�ւ�Q��b�^Ko
oJ(<tP��5&���x��s�R�������h��+�h˷e�~��.�Kart-E2�:$A���t>i[����hg�QjtR�>dP�H�I��������e�7y�y9�,Dy����M��Hqd��{tn�M�y%po��a�|i��$F�p�{ � �F܏_�
��i�h��8�&�8 �u��5l�<��eSMAt�	��n��r�7�U�zS*��� ��L�����v�2��F�l��0�+�H��=��E�Q�2�^+72D�k�Y�]���7�1<�x���z���N245����ʒٻc ��۲m�q
��+� (B�e��-Xdd�e�#x'����W}�o����@�Ql�����<�!��f��}~dh��Zn��Y<t9m��(�f�ll���5>*�u 	���k۰YIN��3Y���Ҭe��6�d��F���j>�:�6�K=*�y���=_P�@">gCG�ǎ}KL��K���!~J����*�6�K�s\��ɑ/wd�::9��,K2֫f6a�rE=��J��8*�N�tP�5<8��\Bw��ϭ�s���;\�a�N�_�&�i�Tl�Ep1=�*-F���Y��}�Z΅���g0��އ��r�X���-\��k�N!<�`|&�ܦk��i�ޯ�_�1��ʇ������Qu���t��wBӏ6ɉ��
�,���}s;�0�ԣ{���y�<U Rq���j	 b��&�F}������N	護�M����L���G=�uj��`��9St���p�j��<�@톁�gQU����]�q
��C���޻Q2���d���z���V@�YX��`^`s:�[ �PZyj .�=~^D�V�<e�z@Z��
�o#�ӓ�|N��v���Wo�5r��`q�����O����h����&�m���" �L�B���&:k�j�a�^��G^��h���+���)�Y>h�o!`�����C����xba$*�e���:�)�T�\�s/�r �4 ���K�7�O��V AKwFҗt�Uu�.� v��n���͘�B��`q �/����N�S�u��������Iϰ�k��2���Ns��n"Kz�!��y%�(��Ϸ)��Ǎ�5HK�n@d-�N����p
�ۚj^k�cL�qm�ʪBY|�+.d.���V0� =f����`�Q_c˷!�J��qg�a��<����Aj��z9q厢����Q��I�gz�`B�2�Q�Gs 3�P횂���O~�M`NSV5.���s��7A��R�l��̭?��㘵Wp3UԪ�c�l/3���N�U�;�������1�[���Utt��Б�8#@���"`w	������>�{���
��J��rMv��Sd�q��$��2'P��h���g�7�P�D9 3=w���6�\�6�̌���`��]��eV
�6��>&��g��~��g/ʳ2~�?%�E�U�t.ԅ��g�
�Q��m��!�'��!��������+ϖ�A�L;����^&ȇ��Vh�(_)�<}4���!`��>X�P��XT��,Q�үҙ
Vm-�xRO
�7٭�P厍o�P
��.~�BgM��2_g����Q3x2�n%gW��i�~f���f�_��&�o�Jݮl���X���,�%'a��;c[�ݩ�St�r�eY�t���P�G��1�� -��3��Yjer(0ɴ!��8ћn�⯳H���N�F��N.�.b�.�< 2�q�o`/�0���2��G/�2�1=�)E��+�$2���d|���݃�Q�OX �I�ׄ��.���4���ɹ���g���#"MV3�E�"�QC�!��뀇)|�4�[�q��ϝ�`�{r�~�4њ̠�m�lU )L��u~^��?���i�R�Q��$�P3��YR��1��#��Ũ��G�,M�3a�E.ĳ�5��ɟ�e�%�ވq���f�bG9p���_�qX1���'��!�����9����QVd���5Q��n�\"��� ��!|����
%�
�y��u2�Rzt�Fz�gvɳ�~�l���܁���4rMfHf/Զ�����3�����h�MP�������Ġ`��q	��f3�x�n�����c��k��3id�!�2���e��,�+h=���(w!$g�n�� �����^���a����o?�<M�y���Є�N9]�� z>�0#e�`�^M �癯+�K)Q�b�j�k�<|Ђ�p�L?�
k;#0Bs��Y~�Z/0�ڪ-z��wa G��mY�㒚sH|�{��T��R����Z�Y�	��p���|VN�g(JZ���a��B�K ��RYe���e��9nZd �G#_d\�4�m�fd�ᚠ��pAp�h�)W��=l=\=����X�`P>bn���1TŦʳ���$�<�1
Q��%%u߃�KW�x��M��<:9�9{*ؤ�|S0���ɣ�Z�ѬLX� �˼ȃ��\d�l|��Y�[��;�%M0:Zۑ&@V�9)����dU����h���L��G����%KV���r���+�I)KZ=21ޗ�O�� Tg��� Ɲ9�.4d�R��܊(� �Ml�!~=�L��
9�3-�1��i	��:e"�L���*�=��O3&��+��μj��$�Ϲ?���@��
��dj��[�⁕�̳2'�`[�$ԓ1ik����v�z�P���r��]�~�*� w�Q��=#3�l/j䈨�Y�}]�a+̌
����4J��YX����x>���7�z��8�+��~4LT��hL��8麈
�B,�8E��N�����6c�~�|��w��G��7�,&��D�2�L)j�rϳ��@A��~v8:E��q��tf��jG����Ij`�]$����`W���x�0}�W� �:��^r,��6�	��3�r] ��k�U@7	��7l;�vm �'0/`l��L>!?��K@U?F~�B�����E	K͏��#L�x߯X���,�|[���y���ъ��!����:�N�	o���y��tL��I9e�?�0��éV���{q���C�D�a�,�9񟦓��k;�.���?:�.i�N�)��Kibr<ZfO�N�C|��4�a�Ӝ|[oSu2nh'G��ef�����O�Cs,Z'x	)�D�# ^�h,�>�'�P%�/7���A�̀E�q�NJ�>yCn����ZP���|wr&y5"&�O�'R�ų�2�,��Cm�S�e� ��m>�ӳS���g��b��g��x��TT<D�FD
L�{���l}����S�M�O�=�6�-+�������� ��"���`KÂ0��K��f]����CS�C����6�0Z���ݝ��x��lǗ_��/-��q�6�D1��v�e?븖-:��@*+U��A�f�kW�b;����,�>�*��#`����J�	����<~b��r�������+Q)[�ߦ4&��cǦY+�-8����2K�rD{{,�?S�9Jg26���d̼��<�-��8�bng�`οr^��nBQm�@b �a�VJ��^�t��o�꯰� �ǹV�����	}��~��p���r�e��%r�6�|qn �������gr�,�媉-��v\�hQ����Xb
�c'�%K7�6ϸR�8�(%�ꛑ�{	V�@x2V%���	M)������
�(:Ď�������u�6�򶔧J (� �F> �e����aƣ)�*���~R l�i���w�l�v��{�w�*���gy ��~z��{�������0ALV`�Lv�`x{��:X�;���3�@�_�xw��98��ٵUE�@��=/�Uiw��0�!����N�I�IЇ=zK��� �_aC�5��W�$^�Q��	0�m0��(��&höD&�}�� ���t�F6��S<m��I5I\"bau��%o�:��ahR{C,����(�I��6���s� �x�T\������4�h_���9���N;��=ܙ�\<��}3�S1�.���饴IT�:ڣ%�z�T��Rֱ�\�f&�$�T����T\C0����$�*=��Ɵ��r�[�H�A(+��<�g	fg��e��
nN�]���F�� �=�Lϓ�#��r��-�� ����8[?K���]y4�*|_�V-����RU?�~���n�r������D=��'Յ��F�z��E��zq|���"-��3ѳB�6��6�s �t�{�h}�����v�pa5�!�Z�:�k)%�
M>~�n|E�e=�{���i�k���g'Y;�y�0fK[��s�7a-4��&�X��] 'Io���/�¬��(�vذ�:Co�7_F�p�`LكM�Yz�3��ٷ�~c��V_����Q,�۰G0�0�v���,>ŭ{��6,w1��uC��� �s�čf7�<l�_���sT����P��M��Q[m:��Ԛlj�5�bm�X�_�n�p�X WĢ����%����X���#J�����e3+[���^��;�z(?J[��U<=���Z�b����T���RgZ���9atJ���՚��D��@�	��n���F�d��������9-J9y����ܸYnW-iu\�[�>n�,�e/����y�=&˪��{���=.7��$��kXj�M���5BB����ъ�]��T�|�">�1�ڏ�3 ۱FF0�	��>��K���Z�W]�LQ%nUZ���f��*���v�r_�P-X���������m^��]饵D��sP[�E�ds7!��T\��4�$0�f9�x=�x�.u%����/�}~A��g�u����&8�[x�Q�eBV�-��-'Ֆ
�+�s�3s�<���}\���T�g8�P��,(��w�oZ�������^����#�?����)H01����W���$��َ�m�x��
�Ė�!���:��D#�a7��M�κ6����Պg-c80L;Fȑ�����Z�/�Ψ��[©U��v�r'1�S�VZ�ۉ��ℬ��.^e8W��W�yR�[j��WŀL�2��f������`A���5�9o�#�!���6���ɪHl�c|��M��:���������Fs\��p��iw 4������o�+��V�F�E��&�2�����hp������`�
���⺭���ϛ���}�2��w`�Vi�~K����&D��\�=�2{hQ~��]�{gR�0�`�j����z?F����Q���Q�E��I��عq�>k81����,X�8�m����6hߞ���`RSv�R�.�py�]���&�sL�"��߭n�U�����ܵ���4��ҥ��y��+�a,���×��#d���in߆� ,�Ҏv���[��v�6`���/>�i�=���9x��wa�ְX�u����ƥ����ͺ�N����?���x�91o\ƛ�-���9A��Y���8k7�oU�gj��9�9�"l��/�Sضb�6@y���JX����N[J��R�κƨ֩wm}\���K��ݶ@��ە_���w�g^�@�,�eU�]A�~�ȗ��u�� ٩�S9 ���*�� ̕�8a�f�}������\1b).��f��Ϣ#�F��N�+�LVy�	L (�vr+V7a���^0^���g���ˡ��S����V"w�,�����(ע��""$�b�z����W�!XC�axz1��Ma��fI�KHK�X �3~��h��ڧe�2c;�s�f�<��8֓K+�/򼜀��:��ʦS���ށ��1��>�yl�n�=� �x�u�&Lv��Q����\1y�G�!� UY�\��EԮ!'��
�[�ϙ]�}�̴�^�`T\��.�甫�e��4zE2P�T.x�6����:��\cKd�,˩��y׫	��F��o{��i;�r��V=���TK�|�c��|�>`�9u�9r�n8��e�l�j(e1����@.i9�� ��}��r6>n�4���p�n���>����>�1\����%ز�W��+s�g�IS��f*���p�����ȒY0z\O��[�Z)�C|9��c2}�Ƙ��=4S�mM-�u�U���O��?����������9�8o�{zV���/��OuF���p^�c{@I͛�R���n�*�a)x�d�vA�1,J�X��ˏ(!ѢN���*?+�p�4Q��ʝI���O� �Z4�x�A�ŕ�v���9+���,��D�ʂ�bF�����~��G��]�cPC�� ��EjV��;RuB��2�*��e'����Q�E}��M���Z�Yت 3L�]�tI�t������=x]��sv[0�WԳ�XZ��Ms����)�(��[����;��Ly�.�GLv��h\HW�SE)�ƩV����9����@k림P���yS��ӫ���R@���*��nx��r}�(��M��(��] 1���Z(�M�����t*� x����a,Y�V�@��O�P	8��O-�{S�Y�YHM�8�O��d���ijb�D�,�p�,43�XDG�f�.-�1����A�X���	�L˔�jف"(�"�"_�y�<x�0XH�����t��&t���� �CaE`����;�|�n>�[>��aJm/^�)�M�z���Y��,i���9d�Yֻ�</]�mGgUN�=�Qz<��a7�"�N���t��п�2�&I��@'/�Nk�����}��Z9��^W�Wx�6nh�����7�LG�GQ���`�O'����v3�;u����\[s��J�^5����v���VK�d�X�m���R����p/w�<��8��{��h��*���0+-c�"iL�!���<�B#"�(u�D�*�w�Y��9CFD�RGi�*�z���x���6l-Y�z�Ӵ'�w-���i#�V���ŋS�:N�脘7&)=�Ph>��=.�e%�P۔�3Yy-��cH0��'�S�=/C�,CW(˱d�K��9b���5hFj)7U����k�S�;��9·{�=�:!�b����s�3X�����=/#S�����2�\D�ѫP���Y�U��ң~I ����S�1l޷��:B#�5�~�g*
2N0s��8��?��4��jf4|4���[=�?�T{���@5�7�K�� �*d��W���ۯe��ҎSY.��RL�Ͽ������I�P�u��(#_b 3[��^�m涅�>~o�j��_�+�~�B�����+�ڀ ,"e�aI���CgM�D���,b^�6�����	��pF���q0(,������`g��e{���N�m�
~�b����"i��z����aF���g�q��h����.hGI%�F�|4�R��.hC�4Ǆ+�/}+[�ְ0�2AN�j�Ş�@9y\}��Y>�~O��2ڨ+	�Tt}�7_%B2A%����%�h��9��nu��؜.J_�O��:��&q|�.�|��EtFG��g��8��i�A���5�sr䚞b�?s�b�\�0��^!�� ֠�����4��9�Ep(�U�[��"N%���%DýhH�i����qB�Ekc�G���}N�?���i]�*�Y�u>����g�I��9������A��){J���p����r����1�f�G�k�rT�E��PI&�Y�2.������l��X:����Z��뿉4uw�G,�j��ЯІ=5�2J,���UP[T�H����<���o��n��ծ^@Oa%ڰ]T�a��yN�8����)paX̫�@��8 ! ��.,f�-@7u��+�u�?�v@!b J�쾷�c� �q�掰Bg������<��sg��;�5l�|�cD��31��Itf�s:�H�Ճ�P��ʦ�y�M�S�F؞o����Q��os���ԕ���q�7ԡeD������H�U��=R����Z�.�������L#�a��_����(�"E�.�Q�t�?Z�_ht�ѥ�	h�)��T��>��'ϧ��I��qI��6>���.~|�هg�c� ]���'��Ka3u�5�ɾ����.3m�0��aSfb��;������o˅���&GdvV�4s�F��F��2fJ���%D��k�`<d�e�-�`p
��#�5�cs8�'����!���J��EX���S�d9Iٵ|�ۍ�l\R]Xd��+� �����] �����sf �¿K�y�"�c4ϱV{���g�k���.���0�¯Ř�����M[>U;%�q��p2kEw��{,��\�m�봣�R��vw��f���Y�Ώ_?�xm@�h$���f^�V�t,�a[(��a�����>!�&k�O �����3Q�l�_�f0�P;	���/	����������{����ɰ0jt������X:�5o&c��l�s�����v�a���C�|�^6�v�0ز �(k�v(� �11�C���1?W�H<�1��g�<���/G]W�9�K��p��j"u���f�f�ٱ�Ġ�EQr���-~��W�]�BbI�͟��cj?�ovǼ�f�*����<�"&�؂;���ێOy@z��$�<��YB����щ��2�
����>㽱�E������o'��ׁ�8>���w�z�>�e&�B�Co��"�1�k�D��v��J���Գ���U�E�so+h)����nO���~�6��-\��Ӊ7��i:Ŧ`_�m�ŵ�)�G�\���f0}	c��� h�t[:��[�J�׽ �u��(ؙuX����� �)������t����D��6�d��9J( h��zx.(�2	/p?��񡺌f�Ur�4v@G-,���e쐳��oPme�r�y��}��Y��}T�ӳ�H��r/�+�.D��)�+xg��� m�� �!�I֥�~ dG� v�օR7:��Q2�X$�ys�	���2�n@�&��u���}�z��Rd��8�$*�u���t�	��n:Oc�(�/`�dh,������쨻y�����v��D}s�
�-����]Y��,{Q2 �MY`�"��k��Y�B�������8������F�����쌀�ғe�{Z�5��R(<�52nf�[��SL���-!� �O4e�ÿY�g�Tx?��WCoh5=4=��g�Ω��C��Ο���m�6�T�X��%��>B�xس�n/�kOa�9Ƶ�8�{<ؐ�K��#ʈΫ�G�%�!I$���@15�t:�����B&�f�MݏS�_� ������s��j��F@e���U���rv{=!X�4ϟk��D�Y��ve?
�Q���9g��*1?{��<�r�B^��!uB��z(��J$-<89JΓ2���A)�ih�������m��`��������)�s�z� sIV����?~W�Ar�}ƤH�@b��d`�@�fVһ����Z��9f{g�	�n�][2u������6L�f�d���(ç���q�2��i��mT���:u�t�`.4Z�]V��S� ̱���ó�r����=(c����<`]^�~�C��<�2qmn�_d�B��s¶}��+��@��тx�Qsm������/~ΎGbA'���Q�xDɡ�lk�,v9�6J_Ͱ7c�濻Iw��Nd��	�a�����/�I�V����[g�^�Cg�ɳG���6���1|�������Q:��մ9j�J'.��:�_��
b�Sxms.E�������	�#G���ۡ����O�w�}v����r�}Y��ʤw���ￃ����Ejnv�8�gxלbIn|��-�ll�Lb �`�G�r��4`)�����s��lz���)X���4�%�Վ��ж<A�ۅ��GG��g�hN�]� �S<,�,P�����lbk���L�C��X>Ň�77oEd�k�:�F4@F�l0�XA ���ާ�N�n�FF~� nT�Ts���"��J�+�u�EdF�������J����0{��7\�2�p_�ν�j�x�O���`;%!KCZHL�5T	�iA�~��4�� T��-�.Ҳ�Ƣ6A���+_�կ�.?�Ái�Z�6p��CD��s�e"-�����|��������ч�}��v��}VàN6�c-:DQ�26g.�jH�"+c�q]�h��@!�]0S�wˎld��d����6�F��['*��
]�2�K+�T�pH��1�� g/�H������>F�H�@� 8�`:���Z�iW�+r 8�=��JKT<'2@���oѵ�6���D�ق��OU�k���:���`����l䕈n5�"�C���-�;9� \ ɦ������Y*��%;=�����Q�G�n΂�r�\��&��^���;�X�hn����&���	[~����g������XQ�@�Vv�8N��5��u�ö�c�|)s�]/u���3o�LTۃ��H�vsdI�r�h^��,����Ԧ����j���<{ZR��C,����Z�� ���r|�1� ����ʧ�D&���1��� v�	��]�"���&G�l�45�=�E;��йc�3xO����f��$Z'��O01��[�tF��L�]�>=��D�Ϥ�a����4t-4�+X�	(�zڿ5S3��d�����
�_��,ܲY@=:��S6Z��J���o}��	
u�cǊF}9�5�E����K<�(;��~%�E���x�	����H��=��J@�zs���G#���N��}���E�̯6�7��1�F�z��U:0�"s�RGc ��,�L���"���B؈Q��j��6t0c'0>���Ud�kdw\�/Nം��<<��eڟZK��0Y����@�b��z0A� j+�]�N�3?/U����:������[o�	|`�#^~1��(�fv'�*�j�f�5������^�B�C�k(�G㳒�X��^�w��T�a�~+�5��|&晬k�,.�
t;�k`0d���[�s��8e �Fu�^���E�1���5��P�D:9�`��;�D���&��Z,��c��}l��A�h G^߻]�FĞ
��]����qrq����hqI���HF�O�<?;l*� �]��p���e�ϴ�E6mt�e�a�8��l�>��Cz��I<�łW�=�'�e�NA�z)���l����M���6�H�!��m3�$Z��f��g���o������&�m�M�ob��0 F�`w��7c/"�6Ơ�Y#����$2J���8�X�5��d�g���ܫl\������E�_�H���ǎ���y�f��o���h?_v(#ⵞgD_���6	IJ�'�"�n��h���X�� =�^���'���E�ei�0bA�,��hF���.0`�q��sS����9&4�<�2,e2h&�٘�lv8��Y`�s"�tα�$�N�V���U9��jFaK�y�3
��0qDM�a{����~����y�%�> �-:�(�yh�G6��n��@�ͥ�����|(���9R��w�2q|�1�Z���I�^S�����cv��4R�TA�.Z���fyf6�Eط�Uw-ӂF�܋����\��1�UCnA���+��knȞ#&��uщ������}��
�gc��u0N��[� ��#l.�)�ݣ{oIؓ��͂�H�z�f���2C�p�%��ì��+�"T�9�6�E�~YN�����Et9R��-+Ի�15@�����w��	�}_��_Fn88����
ڗet��rZd�$?&�|~��y|�Nڡȉ���X�9� ��p��Ū�8�Y��aD�y���Ȱ���)�v��L��a>^�)�i����0ߚ���TշfTrn��t���4�r����5VC�C��Ǟ���eL�ko^g���z���r���SC��FZ}5�&`��`B^L���������%0�6s�A;a:�ڰb��~�,��{7�Et��'5v��y�C����j0E�'�R'���;���:,S����p�E����z�+�22����H8u6Jr��V[L���n�.<����ȝ��О@�[�'B��v�#����-���ū�M��"C;{�g�_�"��h��:�2���a��G_���@N��t�Ow���� ����јq����[�kDd�yM-+㖡�P��N_U�&=��h�Vxoد��`	]8�9�}��3Si�w8�d`�
H9�u��u |�������{�K5�kx�q�l�ޣ=����	c���zo-1.���E셍�⺌���������b2)&��|�	�:cj)Yخ ���fSdKE�;��et[����S���r�7�$�F[�����`d|���xu�nK�̓	�}���N�`	3_� ?�W>)1oek�ڿ|�ngt_���	�\�3���G��&���h�,���3u~�]�R#O�e���mɭ�yK=�Q�����g�]��y@���4��ޔ���D'�N� �8y^��X�^�X��2�7��i��>����:b�����e��-��T����,��o	n&�,N`�J^h��t�����4T�������G��"}#?<�\��e��6��+���, �cN=L��F�5��ٕ�����1�캸��\���pn���t9-�1ԒƳJE��1�� я_?�xm@�|�*�����I�݉�1KO!gDw�z=0J�9*�T�bM����5�8b���8B7YLYkYwv��_�*�F|�^%
W��7[S-d~�=�}1�'fAҎ0}0r,:�%��u;V�E��������n~%ĝ���5Z�-�	���-oh�N��"%
��ZЛ`��"���)�գA��(��Ր����9�X��Ass����H+R��g�L�̀#59m�`OR��|w)����r_f[>bg��U$��9��9���D�,��!�蠌q'i��>�?y/�L?Ј����G�_�vN��4L���UD�ㄤV6ɸ��x���!�l���d�Im���4I��읇�Xd�Ѣ=s�i��M�h��6;R���7�q*]y�z������EPa� ��Ϯ���2�����GswӃ����� �Ը~ޤ%:��`��b�8Ȣ�u�Rdę���.�������5��~+".���Y��4��l�������
tRG3է[7�@@���"�%�8�D����(��P�	\�`
޾��H'�"���a�z��� K�v��L�����mL�9�N����[g=�;��ކ���Y��mF��&%����"bXv��l;H6\�'K;������fҥ��Ri]�����)l\4;M����R�����%פ�g;��N �3�&)��b�x��]���q$��`y�Y�2��ƹZ$p��$��x�MW�)c��q��V��s�j7u�������	��A���q%*���f &c}w��g���߮���`)��p�\�<�M�	� Gn��2�[�tӨP�ʨq�Ҏ�l��dN�_�<�n6����8{H U��ۂZ�c��m�����/��I����&�Lsa��s��5a7��ʒ��� ܚz�9�`��"R���u{�͎�ף�,�K�wF_�q1��gJ9��p6�W{����>��������
��\#�i��kۼ���Հ�4���
�U�E��Q������-������ ���!69~;�Е�`�G��d���8J�,�5ܶ�V�=~��l�h¯�ǯ�
�6 �����ÇO�.k��$2�-N�B�S���"�͟�(��1Vc7 ���(4�n���d�o:YX$��� <r,HR�y��4�eβ�u��a�w���^]����@�&Ǥ$b�h�����V��
��6����	�3,B��ݹC�,��t�ښ�1p��!�6ܔ����]m��'�ĲAc�c����RFY�̌:�{��(M�u@b��.�{u9J7+��CgYG-yhd��ӡ�o���eiKwi�;���};��>￝z�.�6��Ĳ�4J�����k3�}��d��K�۶͌�vp���r��_����k�5A�X��ǟ'q��M���<C+u�s�Dǣ7�9J�����k�ڻ?�e5�M��\�]z��y�0���H���q�"�q�=,��de�҂��ܑ�����pHh�8�:K�����g��{ǽ��t�*��I�N)��{#P� J޷Z�w}F��z�ۀCqoщv���W���<ct�qd��H��3�����?��pz�|QdA�yi4��R�p7N�t�!Z>�,�.�:�^t
�`���F�l��XD*v�n�z�=L�9��s����?ٽ�{ �j�IkOh�a����u0h���%��'�'�b�ݜ�	��X�޽�.�,Q!d�Yb[!�1kK�����F������C�z=f�,����ΰf8jȧk8�{�waTFn�O/x�F��C �>����Jw���4�% ?k[�5s����X�hkgp��=2 S�Zז����Hl�l-sO� e��F�v�5sME�v����L�S�> X7/v�y�L���,=�B$А� x�B/3=���Lf��̪L{�6�k0i�c -�Z�X(bA�s�A��#xB��B��7sP%�b�d�E��%G���D�\̟��?�Һ�Y��V�mQH��,�����
�YM6u� �X�����(PЧJ��h ��h^ԛ�����6����9�-զ�%� �|� ��j;����o@�:�q[�t3�]\�Ռ������*���#}����hzjue� ���6�_���"#����^�<���������L�Id��q�Uv0�e���������Ƣ�XE�j������@RzRc�W�D�M @�i'����˝TEY3��i�'`���p0���t� ST`�l@���D@���<�f��8�����!�����i|R�t�wg&m�4&!��2���8(/�Eã���k@a��xİcR�Qî�.�p����.�tI��h񴓰�q�nh���2��Ss3�q��5v�h�*vBK&�s1VaHz����gRek}��G(�6��. V,��Ŗ�Cv��Am��x�&� ����Vk����Y]���l�����ڠ+gO���q���S-m�33)ב�N�o��˴�|��
�]Eۀ�nX�Eέ&���� 4t	M,4=W1,D(��w�ȎM��OXv\�N���j��Zo�}x%�N��рa#��q�>��fP�Az������i}���+g=;�$8�a�J����q�7��:����7N����}���5Փ���u��8(�l�>� ���Ō��ݽ����fJ�jΫ�c�(�m�V��`��g�dO:S���o5���ybt�M�]`w���g��<G�2F��J�O���W��6�¡[o������@�}����-��O�3�9�TC��L<��YNg1�#l�׿��GpJ�;3,.$����{�܃{�V�	p���$�|��dDQv����FLO��f��>�=L��Тı���f���FL 0��lZ\#�q��v�~��
���:���?&(���r��ɇ�/�iX�Q2��uQN�ƪ�έ��s�W�(Y�<54,|,�����hp*;SA��L�&JF �J���(����P���
���	﯑h7�x������I���ϔF��߽2JL�hN�d�zj�7Kd�pdҲ �|P���Ji���q��촯sQ�S�r;o�F?��#���m0��-���s� %���
Q����잵��+z�0d�: 7Z�
�\u��FD�8[o3=�� R��da�
z�kKo�[����f��(P}�3[����eB��9iE`2�Q��J�GuPvz��0�_,c���m����� &5����{����0W����6N�K��l�*^��8���Z�踣������58U�C�ǁ8�����~Z�h�bEpD�?"�
���Z� f�"t6�*�l�+�)�=3>8Ti:�J���c&�t9�S��&�3�JX��Phb���]�^zܖڊR�^W�W�d�kr;�K���gs����`�q��ю���_�,�?nA���;��o��:�P�&f���XYq��@�6��c�G��q�>������pICFm���9��� �]��Ç�d.X��)Mѱ�F���2P�]�H:uq&�`�}�`#��ga.��c����9�nf(�L��Av��/�<W�#�[̉:u�Lh?�\I�o|��Ur*Nn���y=�����/���)�)
�b�c�� [p�2H+ �ԩ����[���C��R����e���eiy��z�Ɵ�I��Cb9I��Q(U;�i���������� c���S�;G|�m��ᣴ��;\�HDm�еW��[jAß�pZ�V�A�o�^:�Μ?l�O�:�=��,��T���~`����7����kjd,=%8T����~TM�'U�o1'Ci�Iu�0�̮x9D��D��~���.=���)�E�7C�u��������47�d���uw��� u��e�Lp����o�����(� ��=�0/������x�I_"���D�)� �,0�0W/�>����D���<����m��[#L���^�z�ս0j�h�����+}��Z-��&��<;�nX��A<�ț3.���<+��;4�q�MX��/K�(�ϖi������Ȝ8���dt�W��h�n)7���/pذ��(υL��ꁞ=�.���-��e�1�����a���a���Uˑ�^V��Y�T�k[!�t\%�RT0=�Ȳ��s�s�o��BY�u�	D�o�����M����ST]��̑�WXrr�Q,-;a'��Y�p-(d���,�o*���(CJS��a����f_�	�r�����衣�F�i)VH��eK5Z�'�Z4�ۥv���E������V���1�&j��������X�����2�+֖�1�^���ր���Ȉ;���X��� T.1��oh� V;e D\�9IL�xZ5��h�C����ۓ��ewULˉ;rJ��~������� ��,��yF�%�emKwT���bܨ�<���ґ�B�I�u)�_*2��w�G��4�Ct�;t:D�1���Q��.0	B�;5��L��Seݛ6#PV��B�C�G�ҕ f����&Y�f�5��ݭ���o8	�c��y�l����6&:�S8��th�?W,˼_�z-v�+�@��TFD �Jz1�Up���U�������g\Z)��`�7�vQu��tX�;I��\$c��:���&چ	�!1����i��TZa�܀at���^�����ڦ����५�ǿ&��L�K��a�i�w�n��E�϶�>�q���0L��D2�"ڭd�W&���t���F�̽ڄ9yJ��v��[���x ��2gr�]#�UX\��y`�W��BAZ��O���FYl�Q��AX}��:�b��˘埐��̎��ɐa P���7�Y��C�@O�	b�J�4J3���s�[����3b#0����bg*�5�"���%�4��l5/2��>;����C7��'��f��pz�� ���W�˜���{t�V����?;h��^"j��xp���Q�]���VgM���L�_t�r��B��z�d4ʫ��4�3f<�{�O�:6<� �o����`�$!��0'�<�����;�T�2^`��U�r���tz�����r�VVg ���5z� �&�^?�'�@Y�@���՗ �I�w�vx��@G�=�%�%��� (Xv�F�A�����`Y��ek�e��*��Z���Dj�va�sհ�͵��ml��j��
��ʎ6 hs�\.�r,p@�lS�P8��_�F)�&�$�w�
T
Y�$��3�K��v��>P�����0,�L��4.�����EG�s�Yp�+���������26H#A�%�=�;5a���h*��bw� ��
}���6vȩ�������H��̰ˢ+4��S����`�8�0���^����q��Mhe�+ &|T���|5K�\˅�&JT�6� [�Dhp�B��62&5��ƐN;6�E�D�ϰl.������f��a�p���7Un�}����i����$A��u�I��G����^+��I-��a�m�^
��07�6�p�F�������]��P
�G:Z{s,��8�Z�����;�mv}�-=�je�R�c��I�IU����v�m�+����SP��8�o��#�P?Њ~'a�H	H���]~�!�3�I\Q�:S��Y !���I]����2�e�ehyKdcta�k3Î�4	�#b��L&|�)�5Il��̎w�)������8@�oE0[�+�6-���Z��(U�K)����?��6�16���ci�:�gO��_�9n�������J#�c�Y�<��A�	����_���ͳ�Σ�yӳ�����4�<�ƾ\�^�âv
� �O[ ��zϤ!2�����n��u�����M���Y؊l���E�z0�����<��Z�4�����PZo�~ӕv�<2���%��0�2�$,�Z�[�NĢj.�:�\�7yΊR�x�,��6F�����Vd�A3�v:�	�~�봳2��3că lY穙�m�	�+BI�r]��c۽�@a������a�YVa�L�֮t�cv܀�-��4���Ӏ�����W�RWy=�▴�b����Z�s�d}��R�;���r���G;�ɪFD�N��"ǦSw }�q�+�0�Yc�8���t�љ�`�YP�@YL���r дI�����z��7�m���H��]=� �$Z�?���{�勞��*�����w!��u������>�(6v�e��?����[<��5&��f�J��e�,dm�]l�� �j盥�|�������$篾�
Fh��-�Y���?cq\�l#�dcv'c|"�TS��E���J�(���}�l�d��6����A�mԃ�NmN�A�IXA�z�(���5eUS�e�
�E�2Z|�f��������Tx~��Ϊ^Cu7va��	�8�;�d�df L�1H�Y�4��Y��@=BX�2��XH�u���MK`q�P䙧�ϔ&�w����U��6ED�ȟ�O��
<e�Q�Sj�j�F�U��c-�y���j9`���Ԩ�0Wpǳ�)�c\���/o�ؠe���^�R��t��/��5���뇻�21�!������9X��R��$c�K��+�S �����9�rzU0��U[ă	%?ۓ�t8��%j�����J�{`��'-}`���v��� (L˲c2��;�h�����Nח���	�%�]w��� vz*��cQ�T#T^٥������3�쭭[l��i��"�.�����;�p�ɬ��bA�����o�����L�( ۟aT��Y�w!��� Ȫ�l�wE�+B�My�o��T�i�dp�����*� �Wt�̲8m�͒�����������6��,��"�a�:�}+v�5t��+:��E ���q��&ps��ncz1ݙ�,��܅��F��k����I��vZqz�{���s�\�#�6�1͍N#�d��ay���7h^�q|�Ӡ�����V���������t���t	 ���	�7�_���g�戛YXVi�V`�t��V�B)fm��Ḙ@� �����s��\h���\�3'x.���V�\x���B�<C�@JOz��(��.��qQ���k��>���P杳[����J|�0Qܝ��Υ���t���?}�� ��J��K�p���1玥�X���X�t�9]��.�_|�X�a�]�?�o%`]��i�w����DՎ	s��Z\���7��:�0�T�7/���g�d�F����7H�O\��sd�1~M�@�Sc�i��dO��A�U����AqLȊX*�t|�_�fa):8W��R�3����u��ݖu0cQfg<��^�>����9h�6a�
_bΈ���
d���zV;rL��|E'��%5�f8vE��E%��ᙰ���,�m���2-�}0@Z:��}4s��U�O� U1� �<��i�P����ut���j�����x��7���ݼ��%#fץ��F�F���]����5*F�:�%�[����(��ږ�$��g5Q�lF�J|Ks�L�k���0:��6�"��y�V��ϟ)�2I�#�l�	�dڼ�ƭ*lV��,+eu�^�Y	#��ϏS@�Cy{ �9�f��eTeʸ���ty?f|��Y�a�yR���q�¨�ǯ�
�V �A�I'�����(+M�ه3vZ
��N.�k�[��B]W(�CKS؂}��_���d�[�~tͰ���*ǖ�?�6e�0:ζ�hF|�\�ɚ`�]��U5�&�.�x�:G�ul�	��b�0!��h���8�d� �
�[�a�11�r��xe���J[Ѵ&�j�V�5'XYT_��О<;B�t�Jt�u�k|�A�w�`��ى��������|Ѵ;!���a.�/�x=�s�������Y��}��CJAt�h�}H߯r��$أ�9ǵ��v��!gh�:z��vV d����a�l��n' IN�� VJ�L�o����џT!��y��6�y��>���UJ�Oo|SukS�}|=�E�z � �!�Z-8;�ε�~�����B�9z����x�2�Q����#�oE�b�)��*
��"���M�ګ><��`�׮0yS��ă�/�ݿG+6�
3����~�_��4CYo���"����v�OM�r���X-�޶�+2m ��?zN��f�<������t�p^��n|�m��?�9κ�w��!�� �}Z��^�e�JZ�����?�C�C!q6��M7ד��v
a�����N'g�y��܌Ya��4��0 9@F3��	�&�k�����aw?�*��.S�����P��7���lBgC���?�<�!4[���}ڪ<�U7�h�9]fh��G+����W�[�!@��۾V�l��yX�i�Q�_�wnj���pL�eۿ��>�3����,;��.c����>J_�� z���
��2+0nf�K��Ƞ�r�^l��0M܍O�{
���-� �P-Q��de��s�O�&�m��|6�hC�z�7�p��G�C� #�����9|�ƙΓ�]���������t���5�G,��-�.������G��ߏ�T0�s�y�Z��2ߛ��4�ȼ�x��jkf�t5jCG�kz汇	;0@]����(m� Bk/��t`�A��s��2`6�έ� suGj�
��|�u��r�4���l�p3�[2�5P5<����߸^6��x��a))�w&札��"�W�û�GD5��U�����v^+����ݝoe;7�SLp��mGerǇ�y��?�t�+,g��h��wC�`�Ip��IS����d�����cWR㱏~�޲W��]#��e���k�4�4�!��8N��9�sH����b�.�?��O���,��@����d95����~���wt<e��@�{�#"]�@f��ψ�v��d�&��U�}]�8-��~Z�[ 8_���[򛉧��JYhFk��Y��n��b��������X�h���A[9�D��3<z��?=�6L��>�-D� �]`}�΅jؐ�7?+��ד�4��5m197���{�z�jAנ���N��;����t��bp;�Y:^x; �@ner1}7��N��~�� �&P�W�Ŗ�j@�p� )�g8ϕt��R+�Xs�&:�J�e�S�����LaA�ɤ�c[���g����S���ٵ�I�/�ܹz*4��xތ�~D�u|�<l�,��i&�<����K{R� 
�s0k���Č�9c�<wmdp5��2{͠��9�v; �=�Q9z��ǝo�Ow�⯣���{��>2�(��9��5�J�������:�W `��F]�t������R� �����m��0��c�]��is�����TY�5�
 ��<����(���YE5"m���x�z;Ac��x�.�C�e%��#;�sl��<�:�yE�g�4\�r%}�F��5@� P�� m�Z]���n�.h�w�c�qi��VxuVaV�|Ps��?��箟�-E����s��F����%+ �};�X�+*l�P�X����Uț�;���K�~(���|�ɕ3�(��%$�b�ma��>�����vk��!��ú�X�~+�őL�H";F��ؠY��^�QYJ�\[;�,G9CǮ���7b�.ۥB����3�����hb�������Sm��Vr�:0L����۷��B�O]�h���}V�S�s\�W��ܖ�� �Str���>ϵ���p�07����,�u:n��pLۜﮢq�L��� �4 ��!���� s~�ٺ )�:��M�?�*/� 6rG����]���bf���+j���.��`J�Ki0Zwr` ����jP�Lz�R���҇F@�d��f�ۆ���u®c�;A)g��\���H�_�=�ۙ �)��H8X�Y!�,�G��h��&�8�*�@9��+��W��0Չw�.�-�v�� ���ɉ	���K ������e],0vme� �H!5���Z��_�~=jE�sgH�ϋ;�c������3�~��)�l��o�I� �Q�'v��'hA/jP���{!��Xp���FE̔3��z62���B��b<:�8�u�(# ,^?��h_�*M;���E\=�.�8�f�,4��fx?�I# X8�F߆WP���&���ߦ����	.);��|�5�$���������Xk �9��w��"��-v�O�
�G�;��`췉v�1ݦ=_p�ևИ�Ş����&t�ib�}s�ע}@�ބ��f薚�Y�$�M\������
�[3��߸�E���	؝���e0$�y�6%vܵ�k�4�' 4ڰ7�e׻
)p������aǣ	�.�ŭ��<�u�'�#v�k��W���|{������گ"����O-�Ԑ��2-�����#38tB�Ǚ7��9���0N���.�����等� C�D�~T��[
��>#C��!�����o�^�@h���"T��"�L6NR�z�e0<:�SZ��ʒ�ڋ�׮�x��_�ud����Yw#��i���D�0��86IɎ������������zlY�����#:*)�1~������EUR���(��*;�n̲���۴�~o��T*���V��+�m�,5��ݚ�fl[?����ڻ��s,�-�Qa��1�~��ٌX�6��6�9�w)����%��l�O�^�&��	U2��l�F�� ���x�	�8^KM��1x�dl�IeY��?���U*�3Q����̹ގF�<z!����l��y���v�6ищ>�l����:��&,�,rϵs�m�ꍢz� ��f\OD��E�ۜ�>�1�%)��X�W��`�j�2-#�,u�ъ�@���S]�]�~ek� 7�1��"��~�+�z������^%���7->��(�i���|V����]!X�S�W8W�	a�be@��ҧ.����:*���$��Zf`�4�P�s���8pl�7g��6:3Ld�������{�t�<��;���;q�H�����^���z'u'��
cG����!8]��������}��G'(�Aj)�,�Jl�̔�sj�(���+�B?��^&����ٓ��cYA�<�Cs���"4�����s��y�[-�˲�@�LCǹav~�@ho�"��Xk�&�//,�W80k,�{��	��s���@]'!�vZ1a7��i�\�L��2^>]܋W�C7�P6R�z�����K}Z�!��r�e˘��7���r�����n�� Y؝q�͚Bv�Y���$G2mNx/)�h���Y{��^G֨���U<g��Sb~��OM��5dQ�]x�H6��8����A��|rU�=�����. �I7��;��5j��M�q��o��);.���j��. ����$�� ���s��P�H��4#̎]=�{�N���aZ��J��.�/�����iiv��Z	�L����:��eܻu�]�=)uJT�zF���ᮋ�"���7��:��и-�.�f�K�����f
MT���e3�����/ �7y�N��7g�7u�BW��3�);�Nɸ���y�r��)��1�w�nhx~�_�o�7xLg�*�;��(M���׊����&=�$���}.X27�?ǝ�\>�!wa]]��r2B#VA����R�?7��ܔ��^��e�;Y|i�Œ�]�++�X"����� ���I��3I�Ʒy^�.����b�s��u��b�Muv�!7@Z_7?՞�,!�l�)��
��*�'K+n��Υ�8��j*��rs������0=��/�F)�YEc��b�@ ��R ��,@:�#O�yB��]��"���|7��A�4٭ų��Ϧ���#�BG�^�U��/˃��{�v�c�bY.X�s&`���L�(�*g��j�C��cV1zU�,��pEԷ�9@������`�1X6�D�=�Ahۃ��5? ��s^��0��]��\�
�0%����,ƺ�@Ȗ�: ��v@H7W�2�م�-c+���n�%�z&�^�n���8�)a�hm<�xg.K29-�e�R���")ߓ<�����NpĠ� 0�<��2&�uX�MZ�-q�P�
����t��E~��J���n�HQ�w� ��VV6��(�Hߞ'R�m���O?M[L*=06k|�*�Ta�F~�]���^$���S���Z�q���q�=C�{�i glu17��Xb����S�=��9�s׮ �"�Q���ko�;Ȯ�yw�,ޓ�;�5�o�x�:Y�7�f��`BՃ��XT��z��<�p���[o���_,5���g�bZ��!@Z��N��>��'�8OA��X�����G:��ѻ�5����U�������EWV%����ie��<q2-�:A���̭��'){��_����zjG�[8� �����e!�sw	�4:�	 �ge�W����m�JϚ��"��2��=^W\0��2��~�������򗀧���-}��M>�v�E<zjq�ޙ��`n��^���A�G��Ηg��w���Xt���}-���y�.��CJlxL' �ZF��p�@�����Tdx�ji���u"4@G0A{t\��@���m65��{���1��MG�[�@2͎X���/d���[���߇N���Hˈ�t*ܭ����TǄ��
�_�Jfo��a��?���nSN|J��Y��!<���7}�~��:.�DS{"�����-�e��E�  �͌s�*,�󉳇��9��z ��T6d�.����X������:��Fq	�+ؼQ�#7Hjc?AH6�Â�6��&�.�a�aE����YTcC,���LTF�h�,�_�}�U^��a��+�of�,��2��6Z֑إ���k����m�Y�D��&��r���lxR[�g>�(1F?aw����|�nI@�����ٍ��	�����3c�<s�TK0�9�'⇶)mqE�azd~��(�" �g����O���e��%��b\�c�P���s}�qFa�M@�%���H��ގ0^��<	L��̱�_�roϒq��o�Z`��O�
Kɂe�j�����%3���(�U�oޡ��ǯ�
�^L�\���%1:-��e;���*�۱�Nb��c4���u��eÁh�[����w�i�?����VIGVh���z;.X�rB����
8[Y�dh�5���{�0̨b�F?��N���QD�����@�K/����b���p��`��"W�~��gi��ǲA��� �f�S��o3	�c�p��c0w�ӌ�}��&����s���%&�˔��ak�?�IX�*v����0:�����Y��1\��T:₨S���k��c�$\��Sx�T)\�R�	����C�\��m��k�Khb�۠#n	a�"l���s�s������,�5������ �Dk#@Y�:?SPx�yy&`�2�Ĥ�h�Kܟ��-ٶ{D{� F#�; ӆt��R�e�� ������h���ñ��h{�E��s[�^.i��@�q����D ��K�O3y��ǹn�c��9��n��mP�ye=�\%G�ӟ�~^3y���c@j�
��%J��9���y�},���-{t R`H�����؍`:e'd��r��X��o�2��I ��dj�'����GS^XJ5 ��t�X- ��@-#F߂�z��h�o!��v�����5���ob�Iw���<�ͅ��F���7U�������}?��&�T'��<]�2T��e���08 :{�.�}Q[���
���?�O���H��_�
vu�t�K��C��&�@|���V��	��s4o��΢���P���j�qUv���cGd��q�I����3�ɲ$�X�s�qU�{ C`��&U]�a�������ܤ�0dm��,�P�r(t�_�|t�{�M��=���N�F�@Q�)��R4%4�?�-�@7k�IR�S8����r�{�:_"�v�$��%  \�m�����O�syf����
�eQ�6q�%+�+�o���[�1=�=7:(���rtE:a�(�ډ�-85MCl8֘�d�,�qvj&6��+�l�A��kp��$a�Ʀ�;�Ƣ)^7��� �{�e�Je�d�eGэ��Ou@e�y��dԂMҿ�D�n��������8o���|˄?~�PW�A�!;ԫu���q*����?>y��3�X`�p�ߣ&`	V�WQa��F��I�א�uĮ>j�e�)���2L�o��:BME��t����^#��]3���`g��de�t��F� s��SOڴ]���jC�)���`�bP
sp���@��0�q#5[i�N��C��;<��'y�q��64���	s 8�Ab�k�l�����99P��5̢h�*m�W/]&t0��Y�QW�l;ba���t�����f?��CBgP����^��;%�n>U��z���J-��	UKPb��ܦ\��ǌ�mJvjD�68`Ċ��B��l�`�B�ЩŶ�(�u��6F���{ϟ<�^�p �J�3�����ɪ�4��b�X%&a��&��4(XkD+t��픣mW]D}� �B�!t(��?3���.8��g`��T_�^�ք`���k�k8%�5%�=4�SG�+�����gh�kS	�4K�q�f�!�P�Ո6j_O�݉S��xk����|}��K��q<�)���O&�(-ݿw'�����*�@�y�|9�K5p9 J֮�� 6�ӷR�I��3�a0 ����qw��h_�M�.��y�&��a���JP�x�gZ��6 �B�0O>㾟�fg���rr�^E	P�k�9k}�q��'��-� ��4��j���g�$���1�}�A�b����Qx�y����_�r�u`#p �Z�xR�#�\��I�_� �23�6t1��Ub˷���m"k�y���vj��w�h�-�kK���̏ݮ �pIv��1�DYv���w��1���cGY@,�!��e������e���@�w��|�s��(��Y�r�4 ���sL���!�����y �p�Q��L ��V��o�l	���0�<�����pa�	��\�pݗ!��0���Y��6�6�s��N�<�v��VW��k�{y��-����ae�<7 �B�c�Ŗn��-9����%g��4�9fכ�Kze���[S;�k\gJ�lʃ��� ����Ø8�
��u��QPޝ9�U1���N&�� ��Te��h��@J�����F[���s�T/V�����j��usv�:=��v�I�	����Ť%�K���(���!��������0�@���	�AグL���7��K׮�o���.��VU�P`Ы�p���UvJ�p��O�H�vG��������2��7�8����2G���/C�"���)�yr��S^Cm�p5È���W6��Bk��+�-s���"����l �Ld�i���}��7�kkk�6t]����'lq� h�ٺ�$ލ���e��sx���x�ʑ�>Gm�`��&-�]=���ͫAb?��׶���ŝ� ��ȕjE���K;���7�.i$����d�����
��)�h.��b��M��oe�a�-�{��2E] ��"�M ��BY[�+W�-�m6d�����N$w����ڎ�~N����+�����B�V���D�`-�S3��װ�Ι>v�oV(�u¬����Φ����{�^�@�^��E�nj�p`�XXLX`�I���w�a�j Q��^��Uo��S��������RO9S�E��<��+�CW.M>�<G��a�`QVy��=Vʶ�`�a}��}3�����dM�?�	P���垺(\���`��͝�|����i�"�t,]��wOr_f�Z�R+�m>�k�]y�J���K���3��M��#E�j�v�� P��r Q7:k �FJ�v�R�e���I��kt>�َ�F�=�X��(�޴s���,�ZL�_T��񺣉�Ôtq��+X��L�p/�a�_�[�&��r�R���b�%�b�V��o��e9�~��q
�5P��V�x��M�X`�f�% �U(���V``��5�	�d|�,���I1GKb��׊�EH���5�*kĬ���u��=����T�#�g����3�X�cc�cy����2- ��H����NG0��oY��.���͵"l�Wvӕ���`Za���ޫl��O�[f<��]�>?���XQD�?~�`W�b�4K�U10[�ݴ6���[bΨ!wY7d�C���FG���c�gI'jሑk��9)\��G�XYY���J}h�.����3Փd���@��B���H)��zj�*ￍ�b@�^G�=���ꐘ�N�r@��(���-9K9�ͷ�J�|�m��6gTp��E+P��!1̋�g0��)Z�.W�7�lg)-�^� fn�T#�0���$!��t���O�l���N�7�e`����lU`m��z�;c�{�-�l ��~�`a��~�	BmF��h�l4&��$�7r<��o�Pr�r��%�W�ZV8��uZ�_~_�F [vB��c�\:���]���׹��\�:�?��U���*�8lO�U���Ӹ��mhK(�0)���s3u/ܖR�I��N����'��x��~��Ň�$J��`��H�_�Sڻ� �`�tH���5R
ke�������f�1x̞�}�:�}7%��s+O���
��Q0����5غ��Π�݁�N\-��>�xx��Z�^�f��y8�|Z���f�pgp��������P ���?����u�����C���5��)�䉀9�.�<u-ğ�lm����B�?C���7�,���h�}x+u_&��,�ёg wX= �"��������bۀ�K�X�0j���V���Pl�x�y�@��~�� �y}��z0mp-vy�e"��	�� a>��l�m���3J^���}�1"8��=�򹑸��̹�3��Q��~��pQ����,�c�M��G`n�x�g�窶�qŵu�;�j`�l��+�W��Z6��Tf���
�Rf JpNǦ��\v3M����p�w7_�,薉��h���T��7�A������&����U���	�2�w�vqA��
�lX��h�. �,��(��� ����|�vei�q"�iވ�}̞d"鈬�\j����߂aOQ�O@��X}����~&��dܚVB��:\!��>W�f�|����G��+�A��x��Z�>�2�s�����_�@vl���rKe��|I�vsy� �2ޠ�A$�s��f�y �t��ү��8�x�t��cFΒ��0����͸yg����	�� �k���Ṥ2[������Yy�x��kK��w+��Z��6�����՘���(��� �QO��.Q���*;恓5�z��λ������'��eO�(�L3�e)m�N3_�]htu��f�Y1O��%:b:�eQʱ�X���y7�=w5�c�����qV�nr��f��2�,]a^E�
?���s�h�S�z'���>y�(D��{=���_�z� jm���o��I�߿�ô��;g�'���=:�$-�'��r.a)��3@�2��K�o���2e?z'��E�(� �m��󆇲H��v�˯#�v�r������>�V��lm����\7��߽��(�q]��e�� -���9����+�>��Y@p;,Q/���DE(�p����
:�'Q�{�	$�q�њ�x���i���|<=�ۯ� ��`�(e/5;C���Q+pԁ��w>HC���|��oɱ���YD��|�eZ��q��� ��e����k���.-{��,�u�T�o�eݢ��o?kM��I�ggo[��A�\�� ���o��s:�[�C�{�q�Cݼ��0�mm���j�~�/�=�����:��y�}J[�� A<��V'}Mm�?��+��,��Ď_�Zk��:2TjUY)J�
(�j�ј���1#�g8�G>�o�#_h��&�g����. %RUjZK�Z]���߷��ٰ!���FDz�WD����_�s�:k��v�x�/=�p�C1`�k�=Ɯ�� �e��Q��)�2&��Q`�Nz�t�e邘G�C�օ@����Ԁ��m^i��j ڇ���"�}?����}�V(��e-\�[�l��n�X�L�Q����؆Af���V�Ig:_�V��V.p�Mj���1�ֶ�4x��3�EY�la����2���:�el��� �����#�i�&��2�2�nG�L@���5if�*���V�
X ^9R�n�L�o��k��TS�~ Og�0�I��pǨk�8Ue��]=�R�D�N�1�d�}�d���-���vj�@"{��z�D�d�k�}./� � 	@��F7V��S���9�ePl_��F�Ğu0��n^g��FGF3��� 3��=�-|(�W����p[�g��f��[S�2A�;a�"^Q���k0�>��3� �Ɉ����Z��q�=r}�2&���Y�W�|�{��fC�}�?4^|�>��̛���|�C݁'�	"`�&m1��H��j�ƌ�/]��M--a*�ɤ��NS`՟��&l��6�.�Qf;��}mU�n�cT��)n�%�ES�V����`oZ	�U�0���Rewd�z�݊�j.T�-��b�3u!��t���w���E�>����d��|�@D\@C��\#�]>FA��5�ht�4�h�#K��م�8s�ݔ��ݺ�}���6��6e-\@����0�����P���n���J�
|>֧7�E�^�-}��.J�\���2��n�!(tS�V�I�+�;�VN��� �j��A'��i�y�Q�6�n���z�at���Ei@�]�B6�u�~UW�Ry�&�v�X�~��F�-zM-[jMi����:�Ce�.ݣ�)�k�l�,̥��&D��\W�mV����Q�Ѫ�*����	.���]p�dC�ȦG'��̀�u ����:4=��C�[��p���ڞ=�:H1 �+�8��^ۇ���-؏;`w����K
bs>��N�6M	(	�댉Ǔ��!:�?m0`��,���&�m�8n�@�'Pb�&�w�u`'�VXN���r����uF*��{�=x0Uܶ��ui�L�lM��%�K�r
��S5�4�OgH�)�ݏ^`Q��؆q�z�b�Ft��Rk7�x��� ���>mxh@�� ��<�C�C�;)�w���,�$���VӤ� h��C-Ǫ�j������:�ד^�6I��|�AS6�@���Yh`[j -����.�Pɶ>������cr���`2�l��=�BoR,�06$3a�(3lr(��L���3����ʳ�e��.j��zL�>f,^�FvUѭ�V@+�qL���Tnƴ��E|Ƃ�V��Eɿ�K e�DY27c�V��6VR0Z8�Sq�֍�5[SwP�������&��
���s2�v4���}�~C���Y�3e�U��P���p�@��,A����2�sM"c���2�e
W�β��; T�Ԝ)�@�Yj0ҪE�g�ux�=�i�\�� ��)��^�iIMU5R����>�\m���J+��QMfZM�g�5{���\���wfM���?�x�@�9��)'��`"tE�a�^̣�c�W?���ԯ��N��=+�S��q2]��E���͢��ԭ��9�_��
�v�p+T#!5N$
��r8�<�o)nw�M�{b�Abrj�UB�����z�H�+l>����Q6@�^#H�iH(e�p2P&�S��~Ew�&��B�۫M���< � Fl�w�{P�M{�����Ev��� �b``Q�	�FJ�:�U@�����Ϧ:�+�TgP>h�%����ݹ�tD>i�r~�E�(�����э,�糾ʽ�J*���)sm@OU��HE\oo:�̹�� �6\֑(C �w	&bG�2��+w�X���7a�@ �DлNO��Z�}t�O'�F����Y�p��!hv�P�xh=�h*�4c���j�]���<�#(���z���CQ֮��0�}��Y�F�,��h[|>K�=��	�唕��`�S�٢/"�zR�S��Z;R/�=��t�>��ۍh6�c�cY�����er#�+u��o�����s��DS�*@b9�e��[��O#@��K����_LU�)p�v���_�U̒6���;Kwiz�=�r�`br��r���'GѾL�L
fs�Ⱦ4D�D�ru�氀�A��3��گA˖�߹x�qR�}�LN8��,��{�v�eka���������T������cJ{���$+��-������k'd7D��f�@�a�.�I��4�-������ܚӶav2���\�l�)F���[���ϸy�-`)�X�f�Y��Z漚�(�0��"��U�f�87j2'��G�h�ifZ�kI���#h��|,�:�/�c��1 ;mX�d�=��f�Զ@#�wq��^������z,�`�(� RF�G�0��:c����)�VX���p?����G&��%��"����'�NH�c�>cIM��\ ��?�9آV|]�f��ƶK��q��ծk��
�.ۃ�"��c�f���n�uH2[\�)x�ʤ���Q��V#ŉ�`�c�^ �8���3���^o�C��
5L�N����US�uoQ�eZv�O9����Ԟ8y0��ݻ�^=W&A&KfʌgL6�d����L������;��� �9�?�9�`��Xଷ44[xܽ��@�KQp��hE�SD��J���.z��M�!J��ɡlw���k_���Ŷ���� �hHȇ.�ؕ�`�Y��A)���/��rtj��#��u��t���.��˘X���
觜�;t�������ﾗ�}���N�k�[u�r�o�2�>1�}S6{�`d
-\�)�c��T��M����9�{���Xh�u���VA��&����2 5�̔�#�yh ݣ�ʣ������[��EUT.��O+@A2�9��8��l��\�E+��F���G�V����\�����w��Ɖ2j��L?%nI�"��}�x-��Hk��@���;��?��`g~�q��qv|��жV���=�?w*�,�0Nܦk����X�C��9�@�TO���G-�Jtm�sC�=� J��U}���E0]Z����a���=�}3�\�@i �U�z�2z�bx]k6@�����)�p�6w��ϼ��􉠡� =�XtA.�Ɵŝ;�Z3�Q��0B4��ЀqbCK<�zز�t�'�փf����%�;h��/~7��9����ϵ�?}4��R�����$�B����`��mK��<Bstb�71=�D��P�?~(�Q�k�§_�1 ʪ���rS�VrMT�-���Q8����mgi�|K�%��W�o:<[�f�:+q</��-,a��<�/]%��\$�s��r��QS/�ff�Y2��Sو�+l,��&#E';��z��
@������:S>nNjh����ƹ֒N���7G50�wI+O��n�EsXfЯj��|5 �Tl�!��\�
�+Q��	�k�I�U�JZY%((��M{.�m���㨅Q�l����¨�
/�..�h���mLU��:c��W�l}O)���٦�Et��-����٪:��1�۬��g2*�P�ʐ8N�yTM�Ε�
�����>
�'D䷟��<`����R6y����ͩ�A���,�cf21kOb_V+�d���rl$8�-
�w�,�@�;��&$�V4ж��`M Ǳm�?t�V���aƂ��Q1F<�����Ӳ�=$M������Є�����n�ޏ�~/��ȿ�[Vr����nξ��n���� B������"�m-_$�H��'��(s�u��׽*1�q��3�3�������'��\n�o>�D	��(du�G-]�yb�@�ǙPj ��X�6@)����]�*is��jI9��ۋA��R-��S /65��.ZY]d�z?�XrL25A��#�Z�l
��标�W1���Uf�����Ǝ��p�f*����vBv2�Q �?�G��t��Vmݭ�����o�feaϵ��O�e_��0)I��6u �q�+���̔���>��s��|�ASO7�1��*)�ir�s�u�O��}��R/BWi�?��v(	���0�3�V�q��,��(��/~�1s�2���짱(�BA�	!�1��Wa7�\���na&�D��Y �mV`K�
Q~�LP�>0�f12n�My[���=s�jbi�:K�'>JcmP��. �l�P��k�6V �h���Up���^ZkLFE��a����a$�e�A6���Wn��BG����� �p�N�ܗ��t��I�';U޳�w�I�-=� �%��6Rec�ci3��{7����{��9�U�xf\�2���3x����L��}H�lU]P�: ۋk��/��,��Sw�,ͧ�ɦԊ/̗�����
�!�x5�����U0	��`� �`�ٝx�|:Ku_)����>������~��ݚ��p  st��k��1��a
��i'P���:}W��m���.M@�����V���Z<��LL���N��7^G
��d��╫iF�w�^gh�� mK�_?�5�`9{��z.M��q5K�:�ƌ��쳧�Fa���;v�UhQ����J����b��y^��k�>G[Hm>0n�p6ة���>[�S��QRM�z�Q��q=
@��	(�5�3m�w�����0��e���(4DZ����ߗ�ڪ�[���@������-A�?[e��$�V%�R4a�9��x��z����D6<��J{�q��l���M�6{od��β{�f� �׫�Wy}�^7z�R��蹟�w �
���l�!k�����j��>����B��a�dgV�ڸ�%k�Y6x��t�^3mY.��� 6���̺ׯ ��H�2�͒���I��;^Y�l/1ӡ��J��n{�M���e�}�"j`s��EJNa���!�ǩə�#˫��
w�g�Y����MG��SU��by��̡P�;H�&��^.�9z%�m��o�3$���/���q���~1���FcC���ȉ�T����z�@�@\�����5AS����˱����3�ޢC�g���f�ŧ�K#���J2�AZ��A�2%���66({ETm/��
��"b�$�����t��S:����=3#[���w�:>��gX�Y�)�Oa���p����%v�2����v�e�#�!ge���۱��I$-������@�c_�@4�t��0�)�1�:�M��\��v���eW�)�K��� �;0 ��q���s$�A��̑U�Vĸ6n�ӕ��Yc��p�KcS�laCH�Բ ��M���i:��3��ܫ�7�,�,6��鶾�؆.�F�u�!+�\�/]f����E��=]����FeVt@� D���*
{�H#:y7�ԅ�<O���WK���=�%�0,�)�r�LVǕ1\%%���j �B�� U*�=�D�@�>R#��\�aL�8.�N!������r��	wʀ�ޣ'Ѥ��z�	#e�.��~�=��L-�̡�[���s�l-Ꮇ��Lk6���_SW�8�4�:���y�Q��g���#�r.s����S�"��S��)Gs�I�f�r�b�x`���UOK�M����m�x��	�~�\rl�>��K�`k���=3e��NF}���V`�RQ��A�t�_Q)�r�[�m���Y͐ژ��	�7�d3V��4i<]|}n:p�>z�X�>8��\{l�l�i�u@�P-� �j�t����a�u|�y��nD ς����1�1�K �& �k���(L���yz�m�Z�@P���]��8�Ø�:<�"�`��b��:�ibG*'Җ^�JPGh
�ص�1��Gwd�m�ڟj��EB��s����E��J]�$r�R؟0KD�%[gK %~(_�����V.
*Y�*el�κR��Y���%��^��`���l��a�hK9�5A^����D�9G�]zQUq�*�M,��wȈ�X֣qSF*<�A5B��аUPiF� L��N��Z�t��^gVp��j/��˴V	������QI�k� e�D�{$�/��%�R�4��t�֠1�m����>Z'����4o�wL�偌S��gi��c�"Y^��^m��V�C}]�u�62��=چ�{#˘�2�iQ�77�Jo�����9�uρ��B�'
��{9���]��fo�D~���$e�2��o�(�ȕ�������䮡��nU���	]��2A�~0Z�j*�,���5o_G�s7#Pq�%S�ʂ�����z1ó�l��:��V�������(����~��w�/���5i�s��qJ��=S;!�<,� y>�}�M��Kׯ_�އ�`��h*���{e�q� ��z�Ee�����K��*�?$�0�m�w5F=t�o��`%eˏ5S+�V�s���0g��l�ơ �LG��{�C�G�e��܋[97V=ʪ3�<��a�>
'�W�{C�lE�
ڗ<B�j�]������L�6�epV�ϊCs\G��"n|�IYY��EY���&1�[z��!��Vk ^�4�E�lu�£�p�.��{PTB��*@iUsݤ�|�}g�S7�.hb�- H�q�F�5j*�ԝ�z�Y�U��E�Un�����3���I�Y�8��YN��r�VH�n���!�ז��5�3��)�A����ì��� �6v���������g���W�O�<��Q�^[�_MY��~��?O�mL҃�R�p�d�����ðl�ΞJ��\jEt���G��,����
�Gj?�< l��s��`�	"xg>*0EP��Z�����(�W�3ɘ���`e$ԊE�K�䔛�Ӊ'�<�>������\l���j
���O�����.�6��I�a��/�>��|��%�E6��-�z-��HW��f����V� �+0Ȼxj	����7N����	o��<�%�t�u��{��A���;��p��OICl0��|hG�i`�D�#(�n��.���V�n�s����eY�?\�yb�Z 5�]���2��/(=�2D���$㽆�v��Y�����%�s�f5z�����[v��}t����������u�nE�U�u����w��DsZ,FIVhy>�I�]�c�*��([�mr�L��d�]Hm-�H�_��<��i��vjب�8VSM���<�*�rb�zm�����O{Q�����iU�W��>+�@�h�ز������7��j ��C�K�UB�&մѴ��f����x�*d�zߩ�
��T�#.��Z�J@f���%�[k�
���e[�ܼ����o�1�'��7a䄛�B�"����dB�T{�,f�P峰 �V��m��qf:Ȃ�©�� F}@�hz��]���ȁe��o�� �o$5�+�s碾�����Հ�)����ad�����.�r�捬����Z{�����b�|��p�B��i�Ę�oeqD�����M���z���T�H��NY@Tώ��� Iy{o���+��gυK�@o�l`�4�#|}�IYh9K`�Ĭ� A�K����:Ѡ�q���JD��a�Z���Ur�ر�ܢѦ�N���� ��mک�XpN���4�<�5v߇x8�B���C�?�O W�w�&��s���{��m�o�{\���Ap�4\���{*_x>zR�j��)_�Hp���͋W0��u��	8Y��ƈm��.L���:|� �,ت�Ek��]�T]�)_"�4g����T�2m;;���"E����V��V8D��67r����>�e��}� 0-s��h9Q��y|| {G���
��꺾��Y���U����g��Ӛ5ʕ�����i��E>=���)G�&��/)K�"��W_`�0N����!\� ��gRK��V|�3W ̏U�*�D{f����*B��C����X�~[��o%��~bw����&�ZI��Q����p
���{�P���7߈4�ڷ�f��jD܆��7� ��r��M	@��)��MY �0n���J���+�,2*��-!��[��O��� �ڮ��x�>���M�5$�d	�=�Q]��z��#s���g� ��VY�m@U�R̂e���^�1o��%Y�nzߴ��mK΍��9��ߊ���Bi���Njv|6фO);���T�(R���ح}��g����t�W�b!�ʴ��ԅ��O�8BNI.�4_�G�<�2��f�2ߊ�������W��QW	#ƛ�u]0f3V�S\iG�^yXӨ�x�w}9��U��衔(7��3��eY8�"�[�NEYD��?3��gY�W�?��b���v���zƼ�kWd1e�n�k�`��W\h���|����I
�?R���[E2��+�#e���w�H���?�麉δ @[Wt�Ύa��7�Ư�(_��@��sw� X��?F �5=Q �5 �q�8�ׂ��
��l��U��A��.��Bf}�c����}
X������)*��i�9H�"�U3��9��u�mU���4��Ǘ;�F A#e��P��s�z��\`eF�(m~�6���L�1*��	��>�w�^z��wқo����u�LDO]�m-a���Ű��bG|ٚ9�AS,M���gv����� ��k2����D'�\��G0���٧b�-k�B��bSɩ�7�E<D��(�2���`:��^�sWIg���-��؉c���F��L�q��h�
�pw`P�nߏ6ޑ�0bv��X��P���+�h�p2��bj�ID�V�V7�+s�b(x�G5W� Ŧ;O4@O��Uw״9r�ڧ�i
�����*e���S'N��k��pT�i߿�}j ����8ؗz۸��+�F����j�<�u����� ��(L��:ǝ^3��V'y�@��kՓ��{����9ޗ�ih�h�{;��=�p}��7 nToq��#��?�����*�A�0�
@�����h�1���x��r���3k��$�h\�>w�xhq]5�s;bm#����_�}�ӏ� ��O�ۅ��y?b\:V; �jz�fR����'��eգLc�橕��S�EVO5����MTs9����{h3�흺H;�ѓ�m�r��� �{ ���N�q���� �?M��Q���c|�MYAI��77�ll���A�B���������c����Ч�y�j��O�.��T6���Fd��X��������+ �e�;Sc�O1����[6a�2�$؅����a�hT����L�#в�_��2k�9�ժ2�(i#��1�59,W�Ul��ʪ�"]�<q�E/0{�f� +����;
Q��l���Z�[Pg�}���7�lL�"b��B|,k��{H�eN������d���\�?_���%uW_F?>Ggh��R��W��b��3�dG0LJ*�[��1�oh����q�A%��3)��d첢{M ">s���n�e}x�{A��T�J��إ����X	�Mፌ�X�,��w)���3�W��ȡf,��Z����d�|ހ��&�E[��q��	D�D$T�;��?d���߀�w��Z��r°=w�P�}Ez, ����l�%��@�ҫ�h�gy,�º"�oe�i-�y&^�	�#�\K	�,��@؅�V�D�%v7���!b�cw�Nw+R󖜻C���S]���K��|��8������v�K���% UCh�� ��s{Fo�:���+�\<\Ȳ4&_# �4��j%p��0ΡA�2�`"���?�(�����y-�nG�������0e��5���R�d9�5��஋^{-4:�$bQY�f;�������{��1��$��:�Ov�	Ʀ��#����.�X����0���!�3�n[j^�A��1��d�r�d&�Br���i0h�W�38K����H� ���9*��a>�M^�,ق���8��/���	 �� =6�T�>,Q^�B~�T�z}p������c�+$4y��:���B�Rʽ+����k���p�zY*�33��¹�޿��6]�	f�<�\C�J%��Z�0��ғ��G���w��"[`}ł������@�n���Ksi���[w�I�Gn�2�:�*����vC��Ʀ\-!��Ͽ�*K+��i�c�O[��UC���I���Jrq�k�:t2ێUE������"=M0�J�&RMO�y1>kƛ����0FM_����#Xx��g`/{�e����ҕ\ ZI��1��Am�
.ǎ�}d��I��:�&9�������rM�V��/ݎ#��/�a,��p�Q0���i�)@ �2�"�����Kl�gX1&�'c7>�������B��1�%��<�x��c���gh-��J({�2T�d=&E���OW���¡���D@��Hjլ�
Tƅi$�g[i�?��V��:�U.�j�H8k���(����,>�� �m0Q�u�����i�h����\_v2m%`����ɳq���yn�{���. h0�&@�yA��R&$�����g�-3u�g�Uu[��v�Y��r�a�hC�bj+X��Y=��{�4�cL��T���G��Y�Xl�����<�i�#K�z�L�#Nֶ�9>Cn�#��VZLs��[]?�Y{�v0�H�q��_.X*��C���͒���mJ&���.r����ǟF������b�rѓeG���}t@�|�F,~����
��Yܚ0�[C�f&���������#u��O��
�L�0�B��PZm��5�����̏?�<v����n�(xsGf��E�cF��k�`Pv	��n�1�Nٿ�*�L,GJ�T�E:e��������O��,����^z��?&�Ƶ��4��s��F�˪�^�fJ[2���	W�5ߥr��TE ;B��`���It&S���_�R�-��d� | �	P���r�&�M|Zp[~���; ��]\���<�x��g˩��n	;҅Bz�l�vK���L�ӤT�c���g�Wd�,���sg�#i��H�����2J�5z�{��Ы��)E�a`�E��n7����B�:1��xWX@��,���n�S�����t��g�9ۥ��1���ȻT�)�m��J���t��ҁs'��h�`�fsT�E7RU�4�<�T�5�Y�>�,�V"6Vc�F����a!�}�l4��E�; �Ϯ�&ŝ�&t�t���C�O޼�.��a��I���9���E�G�.��;�e���azQ�i��[���h�	�He5�����~��'3�ϼ�Y�L�����n���.�TD���o�D��P�݃���Q�l��|��U��$c��35�%�L�"l������ֱ*�b*,\��cY�� R<�y*�j�T��ƞ}��_���h�j�ٳg��&�,�W��j���Ha7���B��X�Q
��j �2aqʜ��ܺ�{��2ث���5���)��4�)���G&>H] ��xNM�w�)���P	@�3<l�`d%�ޗ��M�-+م`!�1<�r�7�<� aL�N�Ɏ��8lPZah�Ke�q����P���/�v_U��*ҭg]�FK\��α�1���n�¬��u�t�K��˱�x�۳�M[������J~&��c3hjG�E{�v��Z�n�O�d�-.t�%��pzj��v�zdy�F�?p�@O5�g
٭Fہ��:�ec�b`n��2���g[�<Xq#+�q��I��*�&�T?U��oh�yk���O��5��FE1�c�v��k <�����R�H_e�qSN K#Vv���\�����T�?#���!ߎa�d��G���H�fٌ�Y�CG� ������]R���ϼ�?�3���_��'^~���h��߄sOr�`�҄�^:���՘�����Lgh�!���foD�ؙ�h_��	"�4kv�f����o8�V��a�eW�ϒ�n�vV��c�ʠ�t���ΰ��ٝx�d��e�1՜����Bb�Y�"nS�Ω��?5����%EZ�9YJ=AZ�>b?�������.^��N�Aq�*�nlA� �/�rZ�~��elM���n۝����d�4c�c*)k m3�&Ь�M1����yv xl�D�L�2Ke�R�}�6H����& �l.���G���t�+Z wg0��ȵ�_x�nk��:�g9����x��i�:)V��t�~�r���EA��u<�X��
�W~��X��@�̾f��/\L3hW��[����8C08p�
ӻn:��Älsߺ��ґ�G���s�����h�X�Hr`�c����\�ް)A~�϶Q�e��.羟��Jmr��/��N��2���w���V���p%T�L]��n�n����( UT\Q�M����3գ{�B�d�l�q�|�{�I�
�G�����j�綖�}H�+�U�8�V�����m������qƣ&t�X �HJ���2R9~�I��\*�F�Us�B�i�a��B{��t��鴄7S%��MRW�>�,�c���� ���6�;D��e,
���V4���rn;){���IAr&M� ;��X@u��w�SC%����?��[���-�^ô��4��\���0��3������`9��'t+9��ׯ]�]z'�혗
�z�?:�/�Ym�G=��\�@�0`,��������69@���CCÜW�^��GV����uJ,R=Y�`3ԩ�n��[���Q3��j�&�1��Ee�O�z��cVg�1>�r8��D� VhV�V�
��5[�r�+�w9-\�>��*e�UZAk��먛K��h�����+���"Z���Qq��ʄy%0��mG�����	?��x�b#m ����� t���f��Y湣N��N��㽒(F:Qv���U�(�ܙ��T���L���]��[�c��dh���Ԑ�iV�,��T��[=�ǒ�<u�d*�:,7ڵ|�����M�*���M�1���k���i��k�������́�,ݚ���wY��e��q#`�^��9������a�����a��,�й^�����I�����q��������o��Xf@�΃]�A�����/�4_�Ɔ~y�CT+�����@�ߒP�f�?�P,��L8���ي��R�,�>�q���9q{�mn��� ���#�G0$ LQ�}��k'��JvJ�_�ІM	�y�tM��[o��^|>��/�,]��H�����z '�:�i��[��A�i!��s��j��Vm�P��D�g	6�o�$�s7��܊�HʸV��ky�?�X�����D��Q�\Y_��"|%(J�Zuu��ը<3�_Ph�yfEg�yH�5ܯ&<3W�3�E�$��o-K6K@3xt��yt�fTX)����`V����?V��-����v�.��z3v
W�e��(�ۅE����}�5K�z���D�=�y�"\���uS�E2�0u��:�)4*�ђ4�vD����r��J�a�l�g]�-p�$
h�H7��h)���Mx�+H����f,����,��kW"�( wѬj�jι^� ��A�����V�W��n��4Q=��PZ�s�y `~l9mѠvd�ݐf{%�Z�S=�}�VZ� X�c	���iG���g;�Q��7 �aT�(�b��%�G\_>Q�h��c����ɧ�J��$�V:�n�T�cL�Дɑ�Q��m�OӨy �4ש������9k�xΡu����^=���������zw�+��u}�YP�o�H�� 5@
��a��;p.Y��כO�Uk	��O)���a�ع&(��b4�R�~�B=�*dv,t(�ꋡ��� ���Hg�e�iY�\A���]���̍�ގEl̃y�#gv{WG��Q!�(LM�����>^��Ϛ)nD%�NZH7�̐�M`��USE^]p ���rc�,kP���
Z�km&;6�[��\�0��e,�x8 FګPQ��g�ilO!B���z���;�4g��1�٪"K	"� �v�� W6@�,'6�� �i�C���^O?��?�X[��h��=�amv3��ˈm�Y��X�O�K�%�b��F-��j˭f�;��\�Gw�`e�W�T�Hq�����8�\f�((��c:,n��1�l�y�����fӞ�����>�'��m��D� �r�%.�6M�b��.*\��XX�J����xQ��d��d�
J7k1�x��
wvt[,�K�E�]�9t�~�=vv7�TCIo?�����a���EНTW7��Э<��-kv���-e,����Yި�����z�30=`ŋ��G掎�4v]ø�����5	����B���4�F|�]��b���:X:A#��=(%�Ppi����m�4�w��$���˫ ?��=�^~1h�nD!V�&��i�ʖ��gN�*��w�\�>Q�Q4�N������}g����15C�U�5�Y0�'ơ�)؁�X ��|����.�@���Zs+����t�cw�*Y�e�6�˴����z���ި�A�tZ� �ג,���HC+��'���i$ۂ۰����D#C#h�н �*�D�P�e+��x6S����r�-5-���Gg�)��q����4�9�P��+CH�e���k����p�+�y�Y ]\w�1a����s����~�{��-�g���?���h�ه�Z\G�\�(�!�Ǫ���a��'� �%�U��ٞ���e<�;���x+YJN���A��*��'p.ᗳe�(��:�e����K�̙n18�f�/Ǭ�� �?節���i'��r�_��x��^�G��z� qw�c,+�TkG���D�{�ژ�r=�x`���綸�H� �ƾU��8�&�m�[ܑ��	@c�7ϩ	���1(<���k ��*�B�h��t�L��6��G꧘�(F�,��0V��;{��RXY�㲥�V&�2�k��u�\���'�*=�0��h��N��U���XQO"8�J,���jK�)��"��*K�	<|.n5Pm���$���p<}�>�hC䊦�����gmFy�=�����`���X�;K ��5�Ȫ���)P��[�*�M
���Q���i�O(��Jї��a(S ������[��=R� fL��&?�U�O�gg՟*~'�I�H@%s\൉R9���"��L�@��a��og��w~�s$\]��߽�g��#R{�O?Ê��<ޟF:����;�;�w h 7�$ ���A�廘�m����!�e��vlY���		����	!CQJ�<�ߺ#�:�:gc��l�,gE��Y���ҵ�Q*��c'�j�tUg'�z���x�ܾ����U5����J~��C3KN��%�JFuL��?5u�ՠ4j^J_�r�;F9�U:�;���я��{���՗���
f$ǎS���V�l1_ v�4����^��#�ʢ���B��}3h	��N��\�{Ĵ7>���-T�>���"�>ҽ/u ���¢��x�H��{��R�w�^{��#i6��뷯GC�:>����'� �B[���4"j�m�NM ���倽e��#J���~�j���Ik0��bV�����ٱQd1h0��Y�=u����6b�����_�-��4Ap����*4�;u��)��BœA@M�8iʇ�;>+�B`��c��s]��9��t�3 /�=����� �v�)��1P�A1#ZEƣ6���|+B�Ft-<�`�N��Z����Y �j�����!�GI�(���M��J�ۻja#��%X��V�`y��j���v ��HW��e<�`��s��O���<�����z
�S��4�f�ݦ�
�;�� w���`����R�u�T��+��ߦ���/e.ؤ�ʵu�i�q����2f�����:����.�ig��Y� �԰�Ǟ�y�
+�n=̍��jD��z��{�d�c�	�����z#�.�}� E��GۺA��m:�{ә�φ��2"�W/���>��M�d�� ��>�fҁv��Gz��R���'O���[pB�(���г=�^HC\'��QN�`�J]�}	TlVvI�dT��3��u��J�R��D��<�Qة�^�R��P��&��PK�B��^�A��E[������������M�f���r�Q�g�����U�N����%� $�aI ���Y
�V��"E�-K�1�F	`\ R�&`��x-��.�R���6��2@tu��r��_�9T��SN�V��r�h��8 .��Y"*��:ѿ	�_@Q�X�I��~�]r0Iᶭ�b��@��^h��{d`��͒���P���0��&�B�޷㼛[I����r�5ʲHزҰ��޴T9�l��Ro)��m�˵䷷�J-AH��7������^��7�'�Un�WAQh�#M`K �Gq}����8k	pˌ�TO����QG�hVU�>vM��E��L�,Z�KѬ��
��u�5'�U�BH�̇+t&��c��D����n�J�i;�Rvs׭��ٕ�BY�*�W|���v�а�ջf��c/�9J�j�eX���n��Aq��'�L�Cv�}����������ϿH�|�Y��釢�@̋ ��:&h�Qfȴ��s��UL���݉�n{�ɈhʨC�ߝ��rߧ�;�w�j� '@ؿ�TNȁ���6�����tv�L?�(�S!10JJ���SOe �M�����v�168c�X-U�XD������aCP�~���l��2D�ʹ�y{�D��}O?�i!�4n,ax �Ȍܺ��
}Q�ʟ���Q���z1v��~����������y��7 ���X,�c�џk��m�_=�Ms�ڭ �Q]���$�G��As羞��E��{�=짍��-ŷ�6�$�eڠ�Tŭ�p�W�Ӣ&���� $���h
,Q1wj�K���/��������	�#2�D����P.���e�WhjP��e�Lq���z��2ɲ�-��sk����>i�	c��$�w�WI�"�.�I��Q�^�������=��Ar�4�LN��X�Z5e)�Cޫ���e�F6U����
�>K�%��X�}2�j�֙_� �U��uwk����42�Jc�{��(�������"�5ቢj�2�;w.Le���y���	xvH+��2������qFk� c�J�u��,�c���|1���&�P�g�Z��k�*������j�	"-8�bm(e�Q�\B��2\�M�>��{y +�� ��6u�C�R���*�`���\F�(�V�X�\V��V�<�R�+i��\���M�늩�����+�]t�w�񧕟����gZ(4A���ڲ7�>z��O�#�h�qh�1�- �`,����T��2��M�|�����;w���4)\����a$�MP�u [�P�"ؐ��9�~A�l�HL�ƌA�
[�bͰ9(��zJE�[6���T/�����j,9׺�2*V�s��0�,�N|���Q�62^@�������l�O�()q|�y������{�����|�^: ��W���1F�TX�
�1@{f�"��²?M��L�K<βq�쯛�>�P�A��ň�R^�)ujj+K�	�IV{��[�gQ[��m3��v�Vw`.ت�M�bw���|W�(.#D�2�-Y9�hI4�]4:��)���ĥ�P҅{��t�@hk��.�k�6�pm�8�6ȾJ㤩���Y���/G����[�� �\�]*\�'X��:.���7҅���s����F��؇��+BH������ -�z��t  R-�N�)�nݡ���)6�;wa8~?�4�4��h+K�D.�Mr� r���,j�t����RʻﱠR��YG��>N���V�����h���U���5�Iʦ,R~-�]�X�ӈng��iw�K<��.۵_��j �h-<�aZ w>���OR~��� :sd�W=2�H�9y��F3ٲyR+mQ��ֻ D����%x��(�M����i���4;S��UǴBy��ja׆5pD��w�n���JC����MK��W�v��Lݎ A֫���רo���^���($�O���צ��@���2 �[ߧo������_�U����S�f*��|��Zz��S9�K����-*o�)� �����h(]��� �� �r��l�:�ՎNl��rQ�C�a�g�R&�]�@� 옭j����
���h��g��ɔ��[�����m�+@rb ��2�̶8V�2�M����g�}-�t���Z����eL�=���^0�J�q�ԕ�W� ��T9j(h������B�M���g���N舧+/`�069�����0�et���ha�@����e�YC�<R/d�NANl�@{}0�V1�(V���ɌO2l0Lk�T ���vI�lh�a�&FsV��в)^{-��?g	}�`ar[�7s~j��2g�<� �,�=V���F���&�=��z*�6����H@Tr�lJ����Vֽ���x����~%4S�l�ς�оȤ�r�KCY�������� K�Ɋ(�.�Z���̴ �CF_AK�M�ʎ�1��+ �*%rg�+>u��P��K��l+
ϞrR�l�<D+য়5��B�;e���Lc� ��	v%���MX���H�:&,��O������܋�]���?���ׇ��B쁜�i����*�,=�hӂ����Rz�{` �'��A�2��؁	�Bh����p�X��1Ƅe0�B5�H�Z9�#��]l�jzɴ��Kxu@�˨��e���H�K˞<VMb�߃��`z�t��{x�X)�.ssSQ��vTeq���I�E�
5��)���݉:9��UPv�>H���S��5�%YJ}�1U>G�I�F���$-�w��x��]�1�XS[
Q{���YQ�ݫl�"j�x�{p�&+�J��ՋC=�����%��nQ�~f��o56�5-05�����hn�bt�1�m��|gJ�8X�@Vݞ`eh{I�N�tm�/��6"j�a�)�Gh�]�4U\���<R]�q�5��/���r�^�J�c�����p�����)���yD�P;��^M��F�.�Y��{�~�J�%���J�a��
�I��	��jf4:��ك[w	�M1��XM�
+N�E4�r�c=w<V��ʝ�*�.�p.@�"p�m:�Ig�es��ʹ>:�����ki�]k@|@�d�[�U��[�E��y�6�N�}��:�`�L��S��N��7�p��k?���8�a�}�*��;��#u����o�H��!���:�jN}'"��g����,t
�-��q��b�0�cC1�}ثZ�h��x�
\��ˠ��7���w�
��c��=XJ,,j����2�v�<���}�f��;7m������k�k��Xy�_k�U�߀g%�mb^3�m��zC��F�� 0�~"w��{��Yш�5d�`_�)�q��0A�r���(VM(T⪿���L?x�x�|�����-,c=c@�������/��.+HTC��%M"O#~)A���5
=��f}jPLIr�R8�[<ae %��� /�%s���T >��͹߮�?�?�`��s���Z��k];BJ)Ea�U�}���h�g�����%���>�DB��Wm�Π+Syˬ���cVD���w�Q�9�	;U��5�㳅��]��x�Rb�]����5x83aC-���a��`c�t�E�����:7ԍ64s-��_,�[DJ����C9�'��&��q����"`�~�������8�L�{��1�~���k���?3���Ʌ(���O���HA	���0�/�:ܰ*b.��\�,������0��k,Ħ�Bd
�Et��@�ΒK�d҈�g$> ur��N�ΤP��ޏ��F�Dvw�pB��s7܏uB�R��*��6J�$�to�L���Ç��u-���#�bI�k��˗  t�~>}�{����'?I��jWa�nݺ����I�SpV´�����~0;v���Y@p�!�@��2=q4�m�j����[�:��ЫvcG�4�}'|dH���>�`(x�ٗqU>N�=������cu�@P�C��j&��P���u܀-��Յ�eꢑ����5���� 4	R���]�Hs����ݥ�|�i8<v������Nv���J���9:q4"�V�HА��A�4�6�5/��E���1�}i�l{�� ����!Y�YU��pU���WQmA�n��
�f�4��k�f�-���9��|�{�{��\*^[��@�a�[�8p/�7��!�a%��}�жt����Wb�WpT�4���C���2x�$��~`v�з�O=g��Gc���{����6�~ �������F��mR��h������O��|�����t���j��`��#�PW֦�[���H�ڟN�+��ɤ 4���Dއ*��>|���sVh��t���~Z��M	����4�������s�<�~����ͺ�L�/�Zu��|�'Xb�}mVgj����J�Jd*�`R`s���<��?޶C��Y�M���;`i=)�O�{�E��nn��� �Z��� �L�!mG���[��m���ݔ^y�t��w^�3^���l�� �2�j���(WB��4��&�qv�Pi�`��,``w�5]�C,�B�^k�R��i�Q�ѱ�m����\lĲ��� �A�{��z�FsU5D��{�*��]�O�#X�Xga{ ��֬�݄;vQO(@�������Ϊ��I��?��`�o���;�`�����7p�j�2�Kw�.eƖ.����ˤp?���(���6 ,:F�"��x;�zk4�Us(���T�ʲ�a�i���������Ӫ�Ǽ��3'ƌ�]���}�gYN嬆�ă�I�������NA�#����+�hE\_��߬V�8F� �����s���?Q ���e��Ut�Г}g (˱�S[դ���'AU�f�DQ�/���<�bN��·��\�9�hn����,� �#rh�l&NX��i� �m1X���h�������*
1mZhR;�2��N�H�`�h�/�Yx��� x<l�~�����~/z^}���ʕ+��OeP���	ƖJ�2��ڝ��-���P�<��PSG����U&��l�x��]T�0��4��2ݡ�|~a)�]�{� 5 9�����n�@ΰ�w�v���oE�c��HZ奥P�+t7�#5r]Str+"�%X���!�!g�> �e%�YDِ��Z��iXř	�� �1����x�0Ϭ�O��J�s�E�R���ӄ>����TAN�n�J��Q�. ����>`�j���&Sa���=	c����'ja���)�G�Ta�,�S��c��g�����dZ�`�P2�F5U���UϽ��Ӂ�o�F�<��Um0��e��k8�{��T��؀������S�����AgE���m9 ]zD����i�=����?�;�yx�*Mb���a��	Е �;�t�%�ZdFv�2���w�u�y��8:�6~��Q�N� ���1��g�����i:m�¥��Y}���P�  ��c�I���&�)���?���H!����t�,[���>n��>���g\�.Zk���[�q�4q��1��A��� D�|�'85@su�� U�ڹE�w}S/��n~�ظ,���$ؙ���b���Bd|	eh_:�u�L�I�=��D�3�fSsBE�X!d���8Ry���{�99��<�i��ڕ���xUlo��m ɺ�7Yj53��d�uj]Mױ���4��"����ʺH�l�K��;��3���u��U��}���9'eʽ��o�!�D������4h ;ZúV�YU��*����ȓ�r˔[����$��*� Y��,ST4�o�rt�%����*��]h��zh�(ʺ�[�g�&�=����8�~��v���f���/~.����0�����uH�Mӈ��z�6�	%��E-�~or"�������Q���N�ܽq��<��Fм�����e{�����"U����oyϿ�q��O�y��,��U�.�<�acG�� A2�q�;dVʪ���N�̊<@�������/�Q4�yP0�=�;<����T/Ͳ��x�����\(�]C�H�q������-�U`��5��IW�y0w��9f�52V������7��gΓnx#���3N��9D��i��
z�A��LgȰ�ٓ	 ���V�q��u��Х�.L
��mq�1xi9���:%�ú0e�5]<��T�������H��B�'��a�r%;?��JH�U�����e�0O�ElK�8E�Q�>���w
,�1뀈��o�lh���`jF@��
�]k���㫤 w�����*��8�����1bm{v�P�~K�(��x^���DҐ��\+�LE��[,���#X�;v0� ֔n�J�!���r-���!�Ӧ)t,���2��y�{?��.�3+8��®=�8���9oP��э��hbCFL�6��>��;�M���K��@������P��{���$)�:İy�o�0W�w�9X�Ƿo�i|�~���KXz�}�U���Z���ɱl�z�����!X����L�*�����cGb��x[���y�D˘�hN�t��7Ȳ�`U�}��ma��A��J`��Z �|��+Wh��ٔ�uՁ��B�+�`��²�C \�E_z��`���w��j�A��6�H�	Sʭ�	˲˰���N�SXD��ۂ	�su�V8��(�H ����}��#w�i��Y	����5
1�%"@�3O(V
�Cc���MkИ�:>�N���xZu4�N�9���)�tZ�2�b�����"���s�������>�i���Ȟ]�f���ba�Ws��5f��jڱ�{SE�R��A���Y)�2�[QYŦ��f��J "�`Ud�h���>z5�++eٷK6.Rc�Rֳ�tO�bTr ۪W��^���h:˚����������/*���<^�ڞ��L0N�Y�R5K~��+���ԝt%�!�^l�!��v��^�����޻,=S�������O��(��bXЩ�afX�"�j��ڬ
0 � H��uI|����OD��_�O���ݾ=���#}�9�E�Z(6�N�!?�-r�F��U֞G��%s���x�~�D� 9ό�S�KK�fn�1Co�H�\7�_R?�> �#t,c1�`'XOp�e�>�.Q��uƎ��C��l�n���.`b��6x�l���Ȥtt7����x��Eד(Xn�m"��p�`Y��D�q� [Pf���"�Q5�4\b�r��ifh����4�E�[b��Ȏ������!ʶY@#�R�1	�bE�T��B����l��(�"d07Hy=�Dq� i����`Y��F��Լ��:��e���S���9~�x*C���e�Um>sl�>n��:n���i�p�V�`��	 զ���>�Q�Y�HV�i ���e�'À�ލ�XЂQ��aH�fUT��!c��&����+ �K�Y���S��F����
���2�4UBʇ�m��JP�[*��!=�{�Pj�y�l��n�V1�"���8,�V�N�B-ϵ�I]��`�&x�w}r�L+&�W�Um��1�I�����x{��EtU�w�G��6�%:���l �0����5��څ^*��HK."\e|ܻv3�44�aZɸf�]�|�@f90�� h�`T
J	Vs��P]���S��ì�z��f�n2LkU��(�OOf��� Y1�7��x�b�P�gp^y�l*l�V\�:&��-n*���F��xȒ�����-7>��S���!@�#=A��U���nl,��O�%��Ee��i�����/siٹ��{j��=�̖MV�(ivH �ZM�uP��>����0�̛q �f�z�`��ӱ�i�Q_Y���R�����#��}�{����A�G�k�[k"$�V$;��kC�������S�"��@7G���{��6�()(!������vmP^nUx�F��h�b6L�`.��jpx��^���/��8z�HE*��rֲ�<����ؽ���:�v�m��{	�`�p�Wo���3�\
�\��dʺ���-�Ui��M����,D�Yu��4��Ѳr5N\s��Y�B��c�im���(�
eL�Ez��Ǭ�z��� (�^e
�l�$c�'f4������i��JAM��
�c� ��#�?���m�U��ke���32�����������q+~@�6wi�+h�8e湞	n�]���4��i�����p�'�%O2`0eMS��Ҝ��ȉ�`D0&���^K���ޫ��n���1�3�j�5��Zxm��<;+[��@*����������u���i�}�D����Ӫ}X��^V)7f��P��x�P14���I,{TM 5 I+��z��������n\����/����������5R���n����QY�����sR�a��~\�e��޽�f��V�4�:E�*�&`}t���vo$Xl�z�h	�4��Oٸ`�
�6L ��`��҆ ������A�k�s6g҃/���K7����ɧ`���Ϡ���t�����bqu����0.���+O��Վ�4�*i� Y�A�x>��jT��l�&�a�p���0�1f���E}�{������MY0�S�#R
|ר��t|���h%�.ImY���Wo� `���Q�����G��@ҞRxƘr�N�h���%��G���W=�������E�.($�N��½���Y����|5�Γ2R\L�a�>1T�Mð][~?��;_�^���9�@~���Jk����TBJo��~R_:��vk�ǿ�/�"Z�(��W�H&��Ke�[�/���&�=�H9��jX���6���3<��P�*'ش�M�H�{<�<���hufa�,e�ƦcL (�i�Ұ�g��PWc�@AH���z�����#W �n�BkV�~�w7���}gs{S�G�O�M;�Ը2N:���Y��海"�V�NH[�#lP&pu�Z�pPH��hƱ��J6i	��tE�-~��'�A0�m���,�\��S��� �ô���Y�+vZ?�;�5 �0���2ί�.Avf���T]�����rq�rA����ٌ0i��ix
�L��(eaBťȵ0K���F<m��m�����[ aՔ�k�!Ɨ8-cg�c��0�k\S-!�T�3��ՂT
P`��k_�:�\-���5f'V���T49G�[�^+���"ɼհ�2~�7�b�~G��������1���K�X��k.[�
���p����	K�G�y�&�Ծ7sd���,����&ZT�)(����ZД�G����S����rx�f) ������
Б�oi��"�'$C�Y��+
�?t����l���_�0�ۦ�I�ݠ\��V�{�g���|��w��APĘoA7��b�����ŉei�L�z�=�6�3�v;��c�G�u�`��ܨ��\�I8�m�K�e���4;�[iD#=A����?�r#
�gSc#hE�H(D���Ϩ��1�d�#ΉEm��NE��[ ���5�� j�=IR$��:MaiӮ�2��+W/�������:�/�W�<��~��ۤKHӔ�߁�h�Q��IG��^�I{�=5B��4�%�	,,Q�|�aH\0��2 9�O*���Tڕ���'w޿��������g�ш��� ,H{:�5]��;�ᧈ��X*i�O�'����ً��� �}T8}�.��f�!�V���p5�J�,����,[,��͑!���)L�/#F�X�|�7�]�$ur��h�=�AW;�� (��"۾�7���Q=CJ����g�")����2K�	��\��ƎtFeej	}�!,W���d�8�Y=׸�?K5�����Sa8O׺�
>�����hbL�zb�JG�4&ȴ�6cQ���*� �֣�V�M/��f*Q*�,�ͅ_��$������y���k����t=�L��z�֔����G��W!N- ��!�9���ʡ���U�s=��}����?E*l���Aݙ�y`�o{w�52n���ѡ,��8�e\Y��d�3�<1�,�h�]�5�����`S����v$�*��E���&����t�̏I��#�8W�D�=���Y:�Z����tԦ��HC+�ݜK��k�L�uZ�\�x�_"R���l�8���LK�����OG����(���k�1"E�lYwA��M�Ҿ��k�����t�~}�<���P�j���f"/�y�ƣ�������\���X���FN�ګ���ix�!�h��ey,�&��3O��G�H���g� �M�E]��a)�=�A�4 T�-م��	�xL�J�iۍ�J.�wS���[۵�(���!��a"e<��͔�6�JeT�a�<8��#��ү�9ln�h��a�\�e�l����3��ϩ��Uڒ3�Mm=���No�Xd��l��:ƞ�����ݺT_"v=���ey��� C�v�p�����.`
���)�kҭ��Z�����b.h� Ȋ4�S��w�]	8�@7��1W�r�_]�_���C����=�D������x�@z�]�g*A3��U����v�涻|V꽳)cd-� Ŗ��b�#ʴD4IsI���
��%�+�dw�
l���'1�AkӁ��7���{��w�C������E~|�c���}��L���1%�!cdo����И�N��w�!���RP*M�nA��'T���x��bI]����p����_����j�G��̑�;����{Nw���ePLy=�l��.\��+M����!Jf9i^K��-h.Կt�\��<Q�fU�����qw�Hʑ
x���I��}` -�zq�,�ƈ1��Ȕ����⑲D�jp�d:��+�*e�WV*�,���M��K:������򓤘FS�~���I�)�f����W`nja�d��4u�a�m'�_S�	H��I�{e_�2�V��l��7�`h8�zh�Ix8z9J�CS��S7 ����Q�^G
�
}PA����!�����R�@�̑&��\Q�1�Ewiخ6��`�[���A�X���nvh%2������#�	�髟�O:�Q����#��ۿ��	�7��k��Jz���7��ʚ�C;�3�8cm�wQ��X��
��Ԋ\���G��a
�"m5=:>U��d~L��p:�L\T[Rn 1�ʰq%
�3&׻j%f�*�&淾�-ד�]��L�f�35���K��t���+�DU�[~[��0y�6w��5�=��f��նjYov��!$f���=zd ���ݥ�9r��u��<,��M\<o�4�M���Y��V�=��2���"�J��;�uzN��퐞i\��B"Ud��3P!;�a�߿�9LG0w2~C��qL5.�������<�m_�|e=�z�5L	c�.�kk�E��%�.����K#E����U�������i?$�H�	�<7��5b���TP�+��W2�����j��t�,Wz���!���R �~��D[�_��d��A:�\�睷���b3V����g��rv���d��*84d�#ˌCC�	�L��f%:p����h|�2�t�=�7z$5����H����'��o^���<Q ȱ�bHq���0��@��ߎ�$ut����"u����M&�dN�ӱ�#��Q�X���/�&L�IWT�1
&�0�}�����H?=�]y��GHVZM��Ɋ�d&`.�0`��~��ES�
�o�b,����X�xO��)�C����8���ƿ��/�ͦ�;?�]���_~�k*ݐ�j����5�,)�6%``�|Um��1;�O�
�%���B�m�V��±hGtD���je�B�p6d0*��s������>^>ٚ��
��!;�s���쾗H���^x�����;�~�'��|y!���m'�5E	������:��FcE�w*`�Ja2��S�ei�i��؞�T��x}9���z�ԩtPz�
�@%;�@ �B3T��6V�	Z�HM,���K'ϝN\�)ͼiMZ�f��l)�ǰ2GS�2 �ګU�Cb�6�e̘**���9M`c�"Z���B$=�x��&� H��j�rx1-��L�L��=Z�Vv��BD�]5���|k�H8"]�3�Kg��
sf{�.tDe �I��5ꤤv���|߁�� ���;�+S��->���c�q1~w2�R��ب'�Y��X'h��6V\-�F�U��Y-�^O����ȯ��ԝ�9����T=���oG�эשn���ZX7e8~ "��R�|�M� `�4�Mt�9P������G�~�{�x���EjC-��x]y�&�h�,m���
�4�d�M��y�aEJI���P�g��[c(:���[m��3꘸^{����zPi2�%M܀����������f��k��D%�[1�X��(J�Y���������ٮ�Hx�uC�z���:@Bs�2X/�����Q�m�ǒw-Y�<�&FP�'ɂ�Kv��R�כ67���Xp B@�܋�0�������v��:��^��!��x�D�\�ka&;`(�h��t�?)ƭ׮1f9�S�=�HA�!�Zf~�N�ۍ��H��Yx� F�L S4`�|v4����[��i2���u2&w�s}&�VPoo3�h�
���k��f��2��pjGwh*��S��YT�����o���rw�	A@|�;��V���f�mH���mi&Я�g
�y�";w5L.M'.�u�wݭ)��\���dD�F�_�9�$z�<u����h=������F�V?Uw�b�V�lN�����ق z�@jS�r��QRդ/�x�.�I{��!ju�Y�ki�җt����:�����?��4�~_ׁ���_#m�g�Em�,��Srwd�n&)O� ���]�i-�KV̝�2 ��4��r�U�3u!.�V�4pe�V�N����������!o5�wј������nN�1 �����o_��ZOJ=�?�`&�@Z�R�j���>Bae� ]vϾ�V���~�W���H��_"(F�LIz���⩮���)��֖#���n�KM���4]�E�xax:�� t��۴��(�f�#,n괪d�=�<:{i��X�=u��-��*�B�v��k �׮�B���MP��@��ZV�I����\E?���D�:l;�'+of �u\�
��y����/��^���ٙ�^J�ݭ�@��8�s^_��������3G��Ы ������0��E�52X ��w?H7Y����Qk��Z��\봬��@�a���d	c=��1�I�	�GHo6s-��!�N�,�qԆ��� �ȾT!���2?!�Sh�pZ�%Q�;�����h�qw�N\�o�{wn�A�,��4MM�)T]g�u1׎���Y�
���+��0�d�3�����-�ha�X�Y	 �$?��Hs���� Z��>|�I)���o?$]�L��V�l���@/�5Z)����y!4��[��Y�m�hQ�=��cc�'59��x�T����~-�����X�n��i[��y�	�%}Hw��ʦ��ee6�-/���Ӽ|�@=N��k�6
2O�f �)'�H+���\���UckS��)�4�lg��2��
�F0�;x/,Xmj�]ve!&�jC���P���<�v�hrl�F�����71��1<u�Y$�'f_u>�9��Js���F%��z�P���!!�\�3q�@"��qN���kP3j��v�2�wH�[��Q?-w�4���	��pW�MX���'��G;+�d�d���50�>�����7G��݁'
��H�s�h:��;�_�Op鏡������	�?����,R84�T�(�/0٪`�Z���'�]�;-��:�����#lVp)�:J7�˴8O`�c񼉷�ᣂ����\b�s���0L	�J��&�ba�Q+��N-3��� ���6����E��	���~S<�&oq�=�l���oG;���|z0� X�������G#�aj�E� >D�i�)��2GW@m�K��SPdM/��j7��H����X��=2�>���i�;�n�J�O���s���4����/.�k�� �ܡW{S?UM�8�Y܋C� ���*(|��%D�v�?����^R�u�{����ƛH���;�.��.R S��������M����C4��- ]X���v���v?:v��G�^�1���S�m	�*^;�R)<�58��Ho���2�W���t�w�m3&L*׷(OZ�q)���2n˔�?�?X蠷�!����{ڢ�C�3�)��*�1�0n�I�=���$��.��Q���B`<�@#Q�J� �[��Ҩ�9����H#��O��l��n�ISX-,�S��J:c|����V�i�8B�m�Mv�g.$�˓�S�g���w`�CXY8<�8R=դ|M�:�d�D�/�&�
|Vr��#R�E�F�-�<�ڿ��_%�Y������(��@k�4sa޶#��{���,<�1ez1,S�b,����0r�*:{��2�4ud�ViI J`?��a�ԧ&���u��`�� tGO#[��c����5ح]���?�g�Z6 	����s�9(��-�
�hЋ>��Y�`A�14z�Puw����Js�Y��2s+5����M�'���	�KEg�M&p=��+	�@�|d*kV}U��\�+��9����mkb% �b�̀EE�V��t[(���Cg�v_��Q�n�V�	���)�:�͔`xwa:�s�&��9n���E�x�{g���YKY�e�����Uh�*uv6�ɹk I�Yf�����uZzA�����+��
@��4�(k��w�6�IV�EYE�v����{�$S%KFZP�w�M��5�r�;�=e������<Q �	�]z���UL�2)�l�g�8�K[9�������w6��ǅ:���w�^�Y�� M/�a�C���D�75��Qq�*�����:��Y���8B��������8vb,�[t��d����a�\��[���B���)�ޞ>Rm����z4�3��\�ȅ��Es��_|!]%�S@�=�����q\�r�W�D���S&�~���p�Zh��n�J:�bA��0�D7oV
��E`���-����1ЛK7���u�'�j�V���N�Ut6��?��`e6�n��-�*�B�~�8���!��u���x"tV;إz�Fm���� �c����t���Sy��Y��yZ��b=�bV�
;�ȵ�Ը�b�ȯl5P@C3Ԛ��sz���TK��Z/uO��+_}EZ�A lA�
��Y ��*Vos��2X\�>D�oUM�����H	`����l��)3.c&���<���2V*��I.Ue
�M���UƣQܧ�L*��ⅱ�2I�V �~Ľ�T
���BzH�$R��Y�neR���i���T-�#*/�*����������T��Xܞ�T�������x������I�MR2?[�4iYSLΩ&��5��f7n���Z   IDAT�}DO*�j�K�5ٓ-{�3���)����ǡ�����q�;� j���Y!����C�s$ғS'��4���4�u�-���g��ݟ=����ʜJ�m7C�?H���M*�N�k���t�=@���
,7)[��Rz���{!s�Uh�˜�aR�头��\+�|��C�w� ��V����Hwc�.��")Q�mY�]���<R0PRyV��<�_�d�e�VA��]X�6s�ld�2��vX��
�^h�W�Q�k{�7�GN���Ќ����~x�7�pf]<��ķ����s/b����U��+c����{�gǃ�ha�a-�5c!sZp�3.�z�\é�E^`��z�`}��.�,G�2鯸��C�x+*��\����:�n�Pp��C� �Zn^��� �S3V%{L:nb�&�,�@W��U(�������釫)�7_� w��AV+��e�V�ၕ��c�e�ȅ��i����_���x�_��?��		�4��`�sJ�N�q|�gm����݌;����1�[ p4� 8T ,�5Et ��;�Ʊ�}�K����ϔ��Xb{͆%�]�=���4bl�Tt����)��eˍ�7܏�0���AD;���"ҳ���V�k�1��B��&bcA��7��Ke���k�(���Z�`���;*)~n��\�J�Ҷ`e�����َ�-��j����|�g?�k��iU�,�R��é�����e�y��+���,��z-x�xܽ~'����h;?��l�VĔ����T��t����o�y����1N� �6*Lf�]M�c��8���/=���twx(]��xE�̀�Z�_��oc5m)�V�J�d��f �ͱ�B���˸�m��������e;��7��J.����E:�P[��%���"JǌQ�^��:e�%�������H�դ �}�U+�i@�E3�� ����x��%��.�l`��Z�8�Ŕ��ص�c�]�*��&����(l�YL #;�Wp=Ɓ1�dM'M#ߡ[!���T�o 49�K�ʬ�𲎊1MeyV�9gY�n��L�U� u'΍j��5��N��-*���Ck
�������V���~T� ���g�s�iG���v:L��&z�a6���I��]�ᕱ�3���>s���p����M4%����F���e�`a�q�J�5 ��ܨ��W�f�7�'f;ǚ�v$�Z��<�l�.,�^23��6I������^�Z7��0oְјc~�1���D��5��̛Bi��]�5W͡e�]� lz�2����Ŷ�R6	V˙����@�T�V��W�U����(���h
��h �֮���MaW�@�;e�� @뿘��$3�B���YZo�0�u��f����)�L�������< (O�K�ZS���d��������u� �3M-M��l+�wj;k��OF�E*�<?�Ao���x ��kU�@ؙ)n���y�T���\�Bh1c�"7|�F@Hw�
�գf��̾��3���|��܁'
�#�(�߅���`dƉ�g��o�E�㎻~nYf��	��|�����������pYH}]4de�;��u6e�?���+&}u�9�@MKG���e�����o�x���r\�P��1�,���<ܵ��h.�.�M�%��.��X,�Ы�Ƥ��ز���)��E~�c��qA���ʴ� ���d�yk`g����=�aYC9��$/{�4�^n��.��h@�4�~��[1�@*a���M�_淩�!Ŵ+�@kw��h�r��W�st�����Ki��<ml4�A{%��}��t��t�2�;�[T�ё[ߝ��D���s���� �����!f�O��M1�2|�oƮ_��Z��	���&+�~ڇrjz,��J	bC����W����� ��cf �6���	GLy��$�_�V'��������&�9=�0�zK����0��u�-�N�^�x� ���e_Oh����:�� FU��EE�܏��n��ͭt���������
6��aU��<��c�<H}�h��ؾ~�F:z�:�ƔGK���=R`8�s=[0���ԑu�s�d���w��hytE��"�@ڧ������"CA}�
i��3/t!�3��  ���^�!�d����]6�
���E��ѾU2�)��:([d�>s&������S��� ��ALq�b�:<����T�9�M�:V�*D+�>ǹ��y]��F1e8��"j�^]�V���ލ�{���1v�ŷX@�ޞv�����8��:+�m�ȶ�1M�g.�#��H���l'ՃgQ�s@��ik�$i�R��ՍiYq9�1O3㤍qh˓% }TP��h��+��}�Ƒ��qʬ>��0��ϵ%0��h���
M�)27b6��:D��)Ѩ��n�ƙUᬡ�)�-���̦�Cp�y�n��R��FmM��:��kQ��!��Ux]����,�m�����L�ª*��e�A�ŵ��9U��ZX�F�q5��{(8f��Y�f{���s���53P�@P0��fZ9��Ի(��u�.�DBi����y^��M%�z�����}��r�(�b�XdQ(�a�0sm�(���Z��Q`���������&[1��9��4FtR/��:�-�V�������-��+k��n�f�j��>z�K��w�V�`��;~5'�|��X�-;hn��(^��j |4�0��U� d�;����6��ky{�u�2X��[o�Apa����,]��EF�ƢƧZ|K�H��j
F��f��Ϟ[�^�Hs<���G��s�C��6����My�:�8KO �&���ydi���,},z7��O~5�!������.c10�^~�T CԄ 4�$�c�!S`��K{n�y��>=��<�ѿ�$��Sv��T��^���4�C�6�M�09��3@��;��;�hϹH��E�|x��t����O�<���~�."i���<��wRC��;�<�՘�Y~ڎ�,�KTo��[�E<��g�{Ct��-�̳i�[eR."�u������[i�U�Z���s�#6V͓h�h���B�������Z��H�ms��^x �/������󯥞���֥�i�&�U�����%�;�/�_sT�YE�S�g�7�f�3�����m�����g0�xu����Y40Ϙ�@d-s(�o��eͰ�Ӏǐc]Fi?����ՕNM���w<;n@��~�-Ҹ������ۿh�H~�Q�s��l�T�}R�\�@�(�;Ӂ2=a*�ܝE�c�ք0���%��iTW�v>g̱�F�h�N�<F����. ns��}L2Y?����(l��0�i2��W�LգP��ҵ(Y��6e��4h��=�Lz���H��Ku�s��Ǝ�tM�Ku�]A�g�J�����4�2�����u�G7�g�E$#���V�[K�.X0����1|����dSu����a7�2'* F��s���؆}� f;��eV�'�	3�m��8ޖl�mQ��u����-
p.�:{���k�p�l]��̉(�Ak�8�#�)۸#Km�G�_�]���kl��P���ɪ�-m��pc�^?c�e�B.��6R���	8�,,A\�����8��	�7a��$�Ϊ�r#�WP���m��]���X�fU��7 �=a�ÜZ,<��l�#�b�W�N����Py쉂�mTA��2T�:�M��-2Z�*ҋ.���|5��0]$ݹA �Pi�z/��ӕT�U�lG0Ԣ��F�mI��<�њ��=T�Y��DC�p�6-��H��������a�+@�ۡ�]M3,�)�==�iT�U�K4E��p���:.��c5[�n���z7}��Q��\�_ g���R��:������My�K����j1��YQR�9��Cq�Z��B��8��A���I#ǟa<C�:�U��w��
��{8d���I�-'��u����]� 6�t[Rk�s��D~�����`�'����U#�g�6��O�%�T߼�.N"�U�<"�B9Iǅt?���v@R.u�^`���W���Hw��] �.�Y� 0�ڹ�v�����=zL*��mx�.�e�NIa5q����5�m�go�6)؝��D�Ǳ>��c�a#a0�FfR����r�4\-T�`�g��b��|�硇�v�0V	�*�R��$r��1��Rʆ/"�`�*`�Ԣ �S��X�Z�eT���]a��2��a;,M\���>p6�m%p�z6��6U�-s`�s����ȬNܦT��VƝ}�� $*��2f��%%`��e��"���ֽ�$u|z�(��\0է�������ɹ^ @�^S���sRt<G��*��͕�of�e�~|j�H��	���g���Ul��=iP�pr�l����A�]��(����-"�!���|T���&��I�S]��9Z���*�_�&L+k����i"�3�.��2��y*��s�AC��2��0�
Nd��c�Y��4��2�L\%��+�%MK���:��7jb)��<[H: ճ�km8J���U�*�!�u�WLR/��5��w`��0�%���������2��t�Ҹ:sL�l���z5�Q;.��
X�ok��V��'-�S��ꪕ\�x>�n��Q}��@�Ԟ�cA3k��Ol�b�Y�[|X!V.�a�rm65*��n.>7�5�+���,��,Ase'z__��n���g�)����B�2�4c��b�<��D1A[;ژ�P��$P�Vd��9��ӡ��d������	Ju��*���e��U9Q�Q�μ��a/�v�kfa�F��b��=�~50d��P��`|>O���th�kλ� ��ɧ��(K�M'I˻ 8�g�60�{an4�[���^9L�J&Tg`o�i��i�c� Q�Ң!�W_^L/��R슺ٱ=t$]BT�;�,����x5R"L�S��ǀc �Ձ�#�t��M��Y�0�q�9�Z�Nxm%��N؞��&��k���e�1+cAmG�$���^Jׯ�NW	}]=����
�S�[;{:��M���UD�0ݛ%��ì�����Y���o�Oj� G�`��i`Y�C�@-����R;����g���2쎩��G#YI+:�e��MV���GS- P��m3�PW�\K�P���g��r<�y4;����$Ra5�1����cL�6���qVh?;|��:6�.�~�Н�%���}�jЌ)�m����Uv��1����7�_��܏�Qu������!ڝ��[0 ��w�<}�V ������o�Z8S�gI�ܺr5|�x�V1�d1ڭ��2�f}H��\9�ǎ%�9��Mj{�
o��e��&�V��e3M�:v����Y�M�7���z�1�6�a
��p	v�q��\ D���TT������U�Ӝ�%�?�v�!ӱ���*M����+�?Gk��]�(����2M+�!#�R1yNnfj�:�{~~��
�kl���RCF�F�����+��fֱMĮ,��y�M��d��#�>��a�H�
��/�
TV�yPv+���OY ���矢�zL"�����	���@���>�bz��v%x�p�+��.� _�׍zQ3L�ٴ�c�&��D!��b.��.���0L���o�]p�y(n���J��\c���P	Te�l�bJ�{mF����g	z � ��:���"�eT�E���01�{�L!J�CL�i-�v2> �<Z�26�a���+�}2�>C���m<��W�w �-4EK� Y<�;��Ce�S�ec���pNjv����^���� tM�8o�E��Q������^W�#�؆/�̓`��ZB�@��8:�(�t{�s3��7_�w��A�P� �5��aiL���Q!45��0���������I0e_"���W�Ȃ��n:ϊf�,����Vٕ���~&gl�X�LO̳�.kY�U�&h�p��!t4�QŴ�Bu6H���v�3
T\x���e ���<6	ub[©^Gp'�Z���D�*��
n��j=@h���<l��xU`~;i�E���H��Ԩq����~���-a!' O�g�$�`������*�B���*�t~��>���d0���ML������۫��<O��Lƃ�i���~�4�"�>lzI�<Q9t	�P��M�=��v7��JK'�r*^V�jҳ��f,�7��JS��#x-g׼<S��0���A�,�y�$�h]��`�g3�FR0��i��GC�MMhΝ>����jDq���4�Oq�e�^"a:+�6h�e�8)��ܐ4Z��5t%Q6�R��l#u4?���r�w)`DZ~��Y�;_�N��g��ܹ0��*��X&յ���믦��1	
 �2������8ӛ��e��"�=vI���PO)@@Dsth6>�g AP��Lj�d�V)����dy|���'cJQ�`�1#��LK�����iO?���"�\ G���@UW��RC�9�Z�<y�r���Y��B:ˏ3M+k(K�x���i��4p8U�_�1�pYa\�sMG�0����� i�QL+&o lL�Ė
`�L�*�b�0�9
!6�����'f�g�� C5���ϸي@�}�󞑭G�yX˦t�����i�� �%��em:��� \��/��G8��`<hw����^L���z��Z��it����0����*Xf.�M�n�]ۼW������0|����[��\�,�M�"c�I�2"9+d-�pL��2�4�-�g^I��-f����jLW�<�4c��0���������u����ĸյ��^��r� �p�_�ݴR7��(Iק'�2�Y�2�YF�\��➫�f���X��k�iy}��Z5g��� �U��?۱a����l3�l�+�$ 昏,�N6�����;�D� ���"�����D��@ߕs-6�S����,��qRlZ�H�t���.�ER��-w;����~�|�=���%A!�e�À���..����5��a�p�OS0��uS-��s���C�&�`�4��|�~T��TaѰ�����Үv�G"H�G�{�J�{��Y�b�#i~++���q�}�����t�����}��V��}?�6�>������Ur�n�Sa�I�{�߿����I��e������X�-���w�FM���AWҷ���^��:�\�����+��Ԥ^-U�ٝx��ԏ�s	�߽[@DK+P�B���Ӽrkz%M��*���7X�tcw{U�X�-�Λo� ֦�(O/ÈQ�����E�RꩻT���cv�;��7^�d5]�� HI ����ҫ����X�x0s�*��\W��ˌ�f�K�}��N�M˕��~�ry�`�/j�J ���B� �a�֤������@w��W�zTp�+���w�֍��s�� җ��賣�j����v��Dk��L&�i�>l�O��Kme��p�RSK��<l��z��.�؊� �� A%��󌽟��o���Z $���(A����z�����+~/3X����7#-k;5nῄ��-PT�cуcX�x����n"�߻�jӞV7�,=�JX+��f|4ݗ#q�gG*���"c�[��M��s��s��Wש&\�榠����s����gZ�uX	��c�����_ �u���8RV����a��4��y����ϝJ'N �6�nP�?>���mU`q&���/a|��r���Q@eΆ9��I�m��`�7 �۰�I^�B�ͨ�t7
��X��}C�  �ܣ��Zݏ�f�g�j�c��JVU�Ĩc)5+��������*[pk��2���2n���9�����)Q�7Hcj��F�g�㽩R+\gO��EƝF�!��4>�B�R�r���d .��e2A6����a�� j���+��rnŶٴX`(ƀ����Nءir���	��*4+�H���HUƬ�0{w��j���W.ρ^y�%5��;Ex�1�#�J6�0l�ȷ��@J��Ը��94ܹ��C�:l~���܁'
�O�Դ�S�5[V�`�DT>e�]������45+�k�`�	�^�E��DuLu@���T��I�����r�N"?ؾ2�b��6s�A��YD���,Ե��F�
A�@;��>�X���qU��I�:��e�)G{`��:�U�@d��K�����`���5*��Zh%A
�V�p\\n!�58���?Nw0����~�.�1ݰ?���o��o����Qѩ,�;����~jYې�h.�Pr����+�6���z�p�-����� }~��VRf�5w��V�p��i��Uߜ޻������0��/k�{V�1��VĨ��v�'�D���gϥ#�O`9ˮ�� u��^�G��[���g�t
����-A_$�؁C�~w�H�Y:��>}�4�00U������ :A*n����l��t��g�5�H�"-N�u���ϯ]�}�a�H��)VXuų�Ѫ^�K��M���Q�]+�։'ϝ�-4Gjm��	��9�0~^�O~3�	x�F۔w��R��wD�v�I���wR��u�g�}nRR�SSC�2Eb��}��ۥ�_�'6β��Ege��Q<g��
Ӣ2H�Y5��D>Ra�-$ h�y61�k��6+k�̓s��!���/B��������;�����a���>(�CN����<���ı�\g;�q!D��a�4��9����5D���dƵQE���r���ܷ�`z��?�M���;�۸y$�۫lvb}�?�!`�l,��57�lLQz��sڊ�F��N���Ze�pĘ�1CFĮ�O���8���t��&ˀ���U�*c��=c�ʔӴ��ZFGH���6��`��s&�>>��R�h��m�l�c^��B�O�K2�C�'e�iK�5m�c��b����B���"�h�;'�����W֗��)?p�褖Q�bJ����7��s̹����d*��|�4#~G;� ,��<�t��Xw,��2E>3+��&�H��82e���sk�BU�
�`�t����=?M ��/ n@	���*6��4�c[���4���H���2Ƣ؆������yDEr�˲�u�:�lծ6���W� ��m�`���A���BFR�r[|�:��
�b��q�`-��F�$ �	Ea�?�aS��)�r+��޿�3���ۡ������b��d}=Q !�.^-ۥ���r��� A�Fy����8(��{j"�܆A���	�$v��b��j��"]FY�9�fR=��D�&;_g���쌙oi˝5���l�z��E|^FX\��y�qz� �"�ȳ�@�D*��#�.]����	���
�_�4؉v^g*k�c���ֶ����8}�@R�������z�T�Txha�\Ac��/D����?��Eu�;�Z
�$ww-m��� ����H���ɘ�Ap�ß��
dMy	pl �٣��
2 ���'ɀX����N�Z9�5�)�Ɏ��S;�CY���O��O��nþ��������O�z?�\Ks慘������;1���<�N��A�L�-9��|6uU��s4h[����O��F��MZ�7���T����f���hQ�a����O�H�S�����M�_~f��&f���s������?�^z�����~��2;h�tZ�A5�J ���O����?I��h� ��p�&]s���%� �ӻ�=�����S�#���S��J�Z���Gg�=�~�;��n��c���}�Z`wj��-�2��o�͂I�Lr�e�,]��Q�D��#ʮ۰��"�v�=0K�1!�Z@�&���cD�(A�b�g�C��f�^@Zƕ�ۛ��o7!�L���a�dp�7��J�	(�%���i�}�d����$	�(-̻A�����+�`.��̡���(X��\�?[n,Ԭq.���=�Vў8�e:�_���M1���K��>?;x���<����`1�J����q�|�,�2�;S��0��m��M ^�������*<d�*+Cc5?������O�,]�np0<Ϋ��S+���R,�1W7Ja ԷX�A`f�,�n]e<X�%p5�WG�m+�Wv`��bޚ2o���Q��"��m{��e�E��+`��9��("f�C��<�Zq�8�J-BH�~���dZP�$Z��Z�����%�W�=�����xOff�U�鍤��<�Q�d��jMk�?O#MY+�F2�f�j��Íb�cџ	`h_��`/ҁ���Ae�*�ʹ�j�2�c�������b�KjKΙ5�M�E,I�fZ�d�jw8�|����FO����/�	���5Z
s����ؼ���<�ǚ��V����=@���ѫ��4%�+���4�n)������ۤr����6���5���O�{;��S���;���;dz�@�;�pe�DuX��l �F���9y���[A�`��c�S n��A�<�`�	ѥ��ʚ�<LQE-:�4���H��1�c�Yx:l��}�\�w����M��}�..~E����[���tg]i_A�mb�jI��O Y��oٜT���5�	,��Աy�(vE�H��λܬ����r{�Z���i:B�I�"�+7Л�&�0d:����v�m ���*x�Ԉ;Zv���rw���A����c�
Ą/6��Ol�n�,��\�J�����i.�kVޡm2=�����Mu�v�'M�[�U�f�-z#��i,7Ŏ��e�sq�9*���=�JZi=����?x?�Q�r�����Z�������\A���g���`�h����V���{� r���.��r�
�a.l .��کC�8j`+Yʟ�M���o� Ԁm�e�:Iډ��dmEH}�6�1�;#HP֓Ƴ�}%Ak��p���y*�&hO��C�\�T��^�>D�?w�*�lc���洙���,���Z��I�L���4��8��t� �W�X@�犡�};���cA-M���GGf_'P�:|m3��Y��05�^{��{��n߾��<�=�����@�YZwp���Yd|���/a��:=��v�?J��hv%e����k�,�S��C�d���S=�����f��٧m#B��?d<��:C���UK���a^D -�+��d�L1�x�U�/�q"_������2�I/��#��4n�p��4��meq���JؙVX޲*��c�di`Mk������ru�2�u|^��,ֶ�}���*������I*^ �E6z�F��r ��/��F)�Ej��J9�љ頩�`c1�9Q�ϵ{�d�$���C�T�L:kO��WO�io���3mo`�>�	��ྣ�X�4i/��;k��1�f�TW%j佶*��5p$:�(�=;��
�P0΢�*L�����.����6ȟY�g��t|ԕ���력���p�Q'ɻ�N�S��\k���p��+$���t�5u��B ���۩������u�uGm��?�@���HY0�i�dm���+��qnQ����v�:V�������H�����ٮo���#.-�Cy��(�C�?w��lp診'�c:(3�(�X�@'�}EvÁf����h����k�Vy����b�ͣн�Ѯ_G	�C-4^_RV��a��i A����H!�)r�Y���Ï�1A�`�[���[@��f��j=e�%e�A���س��o+�ӗ�t��"fp�5 �`��%c>]@���}/}#d�`��;�����P��Bh�ZvmYn\j��Sb��&3�=7zm ��(bq�]�������r�����Z@k�K��������/�Χ�~γ @�M �+kRK���,���˰b����9�j�M3�(fI��$��4@J]�cؑ+�!ƕL��{a���5 Nz�T����dNwpz�PǦ�ң��E_�M���8Us�*�Iy_ojޏ+w]e��K���|}N��}ϖ#5��j"�Q��O��W�""�O4��oSST�5�H�
��.k� ����Vt����qO������g��|������>��/�<�����{H��"H��_e�^��p]7�&�%|7�UkaՐs�ʠX��}��Mi�*Q_�WU��{U��"~Q<���:�9w�{l�'��a\d�ܽ���	0k�W0C�N�:D*�����*L�-��8�z
+�=i����#|_cG�.�V�VG������]��̣9���'q�>E��B��N�|*���Q�ͳ�M��K���t�x�l9��pM:j���H��"_&��]�V%�Ld<��k�V���2u�ZQ�\��+<�|��iI ��mY]<��Z�i9X;��V������n����K��%t?���V2F�"�"�% �\���ԥk#@q��}���4؇,�{�FC0+�\풮��t_�8n�4��mRkф����Z�N��
(�yn0��-���e�����^h�ܸx���D�ћM�CƌH�s����D+yW�i�Z�L��Ʉ\P!!�ԢZP�ڰ��e�Vݐ���-�z
u��F���.�^c\�%ټ`��m#
��ꋲn�]2aXfZ��M
���h���eM=^ƚel|���Eƴ�}wf (8�H7�eՂ�8m�e7�	�z�@�f�����7N�fK����o�k	�b�Rי�N�l��U�mX1C�s`Ŧ��c�<�G+�������c�n���[��!�,���!��{xt����t���!�r�p�ב���=R R���[J1�+�h��3��%��ag�n��6�N*��p�IK�榾��~7����A ��qU
�.�]]'�h��n_Q��/<&�� ������g�{:��L�P~Y�)�g��,��O����0�$HE�Z�cM��F�,��:!,�ׂ!��]�yԏ4QacP��56�T\��Y���V��!��^TW�}x��i2ZK�I�c��du5��[?�NT�#\^A�s�^iS�E��0
�Va�Z�ݮ�z�V��/>�jIe^���474�!P���c�- ���q|�H�����"���� -���Bg4����g�<�^��_I����5�����0�4��]hso7x��C#�2��e4@-0O��5k�:��4��Լ��g`?(��:�������`�Hi�"���E�i#�Ҧ��qZ�~N0-��� ��j���(���~vu.ƕ,Q�r-��� B�:<��92&��c7z��0'��8�,�b�6�������xߤ��R���~��~����:��G �1R�1f�Y�A�=�G:3�~��_M���`��0^�m0fܠȀZ� �c���Q���:�kS�뤹^)՟mXH�W7�;0��~pc��g���300����}�����:��)����r��v����6a��NK��1Qu�6i!K�� 6y+� �L�%B/!z`��d�Qذ���b��~�%�mD߄vf�jMWgW�bZ)�6�ą������x�}d=xeRu�VI3K�e�	��Η�詨�0�n��1�d+ma$��r#�?���@�u��YHd"]&wbp֕�+5�G�I\�3Z|m���~S�(��N1u9�M�R��Hv^�l������|��:�/.���
榶�� Qn���fe���{�4ؾDF��c�i�)�]
��˞�ܟ�"�+K���Z�=�e�6n	�(f��F9�6��r.ۻ��z�ѹ��񷷫��v� GT�u2&��y-���w��I�k��	P�g +g� � �B�c!���D� �v�%[PwV;,9�����;F�N��1��I8� �d3�*�\PL�A��S�$J/#�b��݄�;;�L�Ι�Mi1[���c�fR���P
��m��<=�>�x-=��1����|i!�����������Y��t�<�>]��h'��WH�8�]��X�}��r��=*��o�����ﾓ�@���n��| L��a�1
���qbj*���2e��G"e�Aj����[G�u�So%��q)x��	�5��wd)X��]{�6��U���wS��w�у�#��j�`�I+-�,���ɴ�XX_�>�F(�]a�V ��k���f���1L�'?'�}.�v|m)��2Ri��X������~�pj�����*�}p�^�����
l��r������J��U*�����V�ԙ
�W*���@��9�5�@'�gx�T��~q!���q� �6n�C�JÔw�Z�u�i��=E������ʗ��{��8�ֺ`x8s8g?��z��t�Z�2ǾJ>_���N�$��;��gcOg����g�mM�3��6�����@5R[,��e��X쪥�ym`G�2����Rnһ2�j{|��V�Y���A�q,� ̴�ږυqO�\e<�+���]�,�?��C�n �����:z�����������p9��
������ڷ��^}�e�9�`���C������|c���(�7��t^8T3n��:�y�c��W��o�����G�.}��'�9*6o�y�._��fa�V��lh9V9����ر��m������\+���k;� k=���R2�h�JCly9ǱhÝ��
��/vl�(�
X���S�R��amһ���h{rY��<�����o�.���y*�u=�8,�*�d�3�*v�bl�3ߴ���	P���,�M�oۜ��k`�<55�h֭����%���e�D�׮Ƶ >��5�︇���
���<�u5�A:PC�J�>�)�3�K�&�s���*6RP���|�0���c�- N_dC���I'�}oJ��a�"��mh�
�r���3�ds�n����0����e���,Z��F��ѭ ���\���f`k�)۠�>��	��s<ƻ��&�����3�����	*��A��CΠ�'�N;K����������"���r��3N~B��(p��F�@!�v1�BH���W�����D�"h�����|�k������$u��W�����^��Z�/P�:���!E���!m�n�uxb� ���;B�A�AFj����G1��έ�B;U+@XP0���R�dJ� >?[���4K��)0W��a�?�4����R?m�o��?���e�6��ǈ���P��+3C�_�2ĉ/��J�KeJ�����	�{̎%��-p�d�p��.�V��ՆFDmN��7��1AR����\w��"����Y�#� �Bٷ�&���_�3�&����_�c�m�ѩ��؝Gv�i+�ߙ#58�n��[J��2lp��0��������1�,���q�y�; P�T�6����hZ�{��JL5�����qƪ���xf:A+��Bi���^B�\����]]O6
�	���V`!����{�h/0��w����㌉�i�ꭕ��H<�*�o+����9�Y]O����Iy>�Đg8�a`8�����1��s3�%5n������ӎ�*�\ķ��JE��ە�:+g�Xb.`5��~�e�jg�~����-��&/�����^���.;���A�`��ׯ�k�g����<�^}�j��ҙj���Ơ�uD�U�W<0�^{�U�|-4���"����XD�gZM ��О��e���� �U����� ��~��L����Hmlf�^����)�޲���b�)��)g����E�h�j�O�,�Ȣ�I�)&SF�*1-A
�ο��w��Z�ؙ��9ÕX�����D�)D�ռ��q$�C
^�v��bӤv�@���B��}�����Y*��/���fx/�񵦨71��X���gz�l$3�c4�Ռ��ӗc-(��=����g�q�����p�B�ꨯ�?�
��-\c�����\�/�- bLԱ&�s?�P�Qb�[I�R2OE��6cvKk���IkF��d��l�+�Ӯ�M+��Ǭ��,����F ���2���9� �ۯ������9;8W���e�u]�o�O����BiEnjkc��\3sD�Y�d������]���P����e`�
��ryk����� $N m�(�D����-r�16��뇿��	�>__��ح�����ĺ���ы&���\ ]T�19k%��^a	�i|� �~��3��$��7�J@��<�gSZVG���(�\)УHa4?�G���1����5#̬��>��u�BĲt��޻C�$�@`ɯ�����/W��4f�����`�6α�r7 K>���ZC<��q�_���{.�����
"*��K�I]�A������{���t��z1KO�=i-+j�6�yŒ�(m&xd�6�{�Dp���f�.>���^IF���;�=7�����f&X��+FH���������t)>�����Rخ��� ^F|N�J3H���������s��_W�Y�����h��P ���Nb�h��w�ҵh�R�{zw(=�|5��l� WQ2OeUE�\�{�]���w>��y}��6̂ӣ����������Q����VE�q�1���f�S�nZPL�����V9L�� ��Ы,�� [��.X����g�W�� J��vE�9�m�jj��3��2���W˱�$
BDL�T_��c�^]+T�x|f�3#mq^�'�1�Txv:V7(ff����E�8�*�������e�N��������=��E��:���t74�&�a������������Ӎ;z=eU^����u�9>t��(*-cG��+_�x1���{�E��?�����<\����{?��1�e�(��<Ev�V�7Y_�S��7�½	�x�F��gu/k���p���3�bU�:�%��q���,`h�۱�u��*L��%E׻��U�|o[� @��l�,㲪�����k��U��������������|�$�C�[5�w���C�D�
Ɛ�G�A�Y���q�nI]��ޖ �ɸ���jj���k@lQ����k6a݌��)��MDJ"ǀ���h����&���MC��%-<H-yX>ύ��H�d}�W��ό-,�zd
��ez��!�P���J�uShl���`]q�����E�qe.7�t�s"��$ $3}jc���\mMݍʊm!{�F~4;��ќ�N�����߈`O����O�0��Rt���
��E�#0R������%O:���^i�@�xM���1��vP6���~0
7̀K�ɨ���f�m;
��BZճ��##�@}���j0S1�.^7��vu��3��Mu�Ė�������$�s1��Eڝ�e���_T8�������AK7���,`�0�S�]�=*gW���gّ?H7���?�K������>�����#���MpS,U����P��7DК�Yf���v�_���*B���H3=T"�-t4EU������.��h%H���Э�i'f\JqW��!'aG�/]#}�>9�Fg�	 ���@#��^�j,���36M��ӧؽVR�})c� +eA���ͤM��K���
��\|e�`��'xn��:L��:�= ���h��KpB��3���セ@;��4���tm��8�憧��ц�`�Q�����v �ZZ$�TM�a"hw��Z�S�����;w.��S0%
�=W�s
0����2F�+Y��b�7#:��^A��3I�"� +@Կc�th>���j/���)�g�9��C�<���?��/���F� �?�Mǫ��?�U��LuB6���!���7�}y͚v�IO�x`V�_�/� b����i�AQ`mq�i����o�qT/�D3׌�I�'��4g�0���w`/҅+?�ǫ?�Ǧ Ӥ��!��
Yq4c0�^G����)���L@`� )!���q��hD�]�L��hL��ښ��@_��0xo
�8��W����+p=���WF���0"��RՉU�ug�R�685e�g�˵�W�*:כ����
<�@�1�ǡ���.c�e_o\H t�/)V,��#�W�(�<���!��j�������E������ӥhg�V��J
*(t!���i�V�Ds�h�*��3}�z�FP��P%`�8��n�/m�\���h�R�g��T����5<�.�s3=[��[�!<�?����]����qT�C5��I�Ԗ�%Z�٫, c�,�i�{���;��|�}ށ'E�.z+%�ASk�n��v&�x0B�Vmd��v���̧buu���U9�>�oLY)�-�����<�$�56�5�х�4�Hꂅߝ��!{��;^dQ`�����ñ?�t=�����/��g���F3���X��t�� fM=���
�Q�2(�- ��� B? ���G�P��iC�0��*�l|:
�!˥>�*�{��A�N�uvtq��(�V�a����^�/G��ح�k�F��Ψ  ��g������XL����l3���s��/�D0@����f�j�,��81�8�Ċj/�ȨYR�Xſ~ �8s/YtF'��l�%�.�6��n����8v�hh�LG4d��>�s)C��F��L��.֖��&U�<�G��CR)+ ����?�zk��)JdaR <�4LaH9��QZ��rײ w��O��v�=�����XZ!0�>�eU0���N��)�x���4N�S����<'*�¥m�ڨu�K
�C��8�j� �@�{�l��|^��0��y������M��x�b��kVΫ��cG��R�jEh�,綝K?"�a�xl1�V���@�¥���+ ��t����y:��]�t%����S@)<�sR�,�J������Nr�!�YL��F�lYRҌ��{�Ap4@֋����*v�^kVZ&�S�/�����#�4O��nJ?{��4�xm3�&��л%+��4���?��),��Q�B�,m��p�����t1`���#�����F�q�H������-��Rh�Ж�b��ݘ�c9�Z2�������.�it�a���Ÿ�����*5+jJ�g�u��v�;���*R��.�g�S�	ᤘ���^0�^���|�iCӃ�|��j��^�:�VR(�0�5����h����h��gUd>Sn��R���J������տ�x-�Ll�bk��-E�K����dV=�y���!;M�en�����Y�� qOB ���3x)�ءO^��@�M����$�)w&u��9�:������	p�.�~�@#��MR��v� � ΄l��w1c��Ea�E��7+�͜I]�`�3�:���YXp-Kw�J�Z�[r���6�<5��l��J��s��X���6�N/FG����Fn���SO��yiy�ŽMZ���O���&��QUFGh]I�s3l�������63��_�t9uREdۆe^��uX(�>�kr��ľ���Ӻ+Ӽ�&>.OS���7ތ *�2�6۰��v����U���A/�2e�n��4��r�\s�����V���O�d� t}�'���b�P/�A�����W^Pv��v�V7�
�4�p�s#�;T;��2I�6�Z��1���&��d��<u�x��E7dٹ)��1�\�4������m���u)v����ｔ�_E�s��v�,��Z-t�%�8?� ����5R~��6��)"Bd^�N�}x(-�>�]5��N�.��(�H��]vح�@[�8�0�#�19g�ܪ =���g�7Sx6wŎ{�N�<f��((m��Ze���r>��#ҠY�_��r�I�x ;� ��>W���o���6Ə��s������!�} K�d�bʀ�#�ˀ�tW4x�z[��9�:q3H�cz�����Չ�1���0�TOǵ��e�1__^����wh\�9L�5�~����ӻ|
t�9Q��וY�Ǭ�B!��8F�� K���:��)�~���ߊ:�⿣HU��S�SWf%&�2��pv�k�:ؾ�D6 p�%��� b�>4)|��O�c?�
G�mnF4K��o������A�j���I�����Ń��2��?����T{�c��oQ㼌�|�`�R|ݯ,;j��f),6]nO.���r���
 ��{�j��m�ƫ�����Ϧ�"
V�Zf�H#�x���W�����#�2�v1��D�K;��pжoQ��eL�c����=�]E����2ť9c��Y�"+���x$8��#ڮ����:�_aɑ��y��H�� �4�w�z�'��O�x�@���E�;�p6�c9�1�M��^|�� �S˄���z;Lw���*�N�ob=u� U��Q��%�ҷ[�A��0DK���A�� �r����I���������H1�a�<p�.��Z$�&�Q+ ��?5�n��.������g���d0� 4=hHnܺͱh���$�쉪��@�����}�i��И;v4��sO�r��޽��u�6ȹ �>�L]Sm�G�a���$e�Ҫ�,�h@�{u5������	��	r�6�>XF7��g7T᥄�gb�`L��ı�Q���IYp��7����Z#ShSXH]u�����S��d�]�Q>GcL�ȼO%<sԕ;�h.!&W��˹���5{:���mz7��}y9Ҁj�|.#<�6��HU���5��Y�i��=SCmT6Bd�[��cWoEߡ�_���u�ꅋi@0K�J�\��fTv�c�������b�.�z��Q�&�#0�ZE������-�26:Z0�E��_��]?�
�����g�3���{����`Q���{��u����-��-���0�D��Ӈ�ү��Wӛ��������^��kj1`�6�j�q"�0]������m��.��g+����, ��x�����q�կU`�`zFpXÜr<.��:s�0F5��������~����|�����
�8=y2B$K��?B<-�"�`P(Y��~���l�	vTƅ?��Y�1���\[�+�lF4n��ʍ�A?ļ��=T�a��\Uڟm֏M*��T[��d�`�m���E�n:�!������eu��>�����殮U�x��<���"��9r��,d d�͊<�ߕ�K+<�QY���d@0��S�R���z�I6q:{T�<�I�$�g-@�X�{[�A���k���3��`��mE�^��"���'_�/�p����jp)���P1���Ƙu���_[ċ�yE�{<�I�:���7s5����d@�=�^f�Z,G?���%�{�����z�(�0��]ޛ,�)V���~qW�C&�U`u��h�'�l�D�����8��=��r��\�� � �%(}a=V ���l�]zs>�RN��x����ewl�e-�ie�+���,%�hC�{�S=;ރ�{��_�9-H�8y*Ġ�C�f� c\٦gi�W*��-��_�p�pЫ�j<�~8����k��X�K��X/��>GK�[�n�s��HS<�?5����9 ڟ�����B�!����cP�ق�"n�׵��T�L��~O�]�?��,�=2He.�2@U-@2�h
�`����NL%i�B�Y鹅���2�:�	=pJ9� ��,�(١5���;q��a�V�q��:�U�U<E�f	���-I��~���Ѳ@+�"�	��Zۗ��MS������]���x�"�v����G��Eқ_��=�c*a��a��Н�J@���ө��m��i��.e��4t4����4x]��ZTqϪ��ԃȊLZ����ˮ�U`�}T�%�9@*M�%響 Svjǔ�ٔ&w6�M&�:����s�����]�elԹP-	��.Xre�-����Cܗ ���:���G�>}�{�2,�M�Ռ��u%਱�x=\��S'+?���>���g�%�¹��p6 Fk���2�3Y�+�nP�F��@%Xwz��9�� a}g9~$�����a���N���)���"�#3�a���f�Ǔ7�F�{1��d�br���"e��6�]�}o��Q,zPI49f���2c���	�t@�Ȕ�D�;�_�ՠ�R���iS�$E�q"�T�%��G6A���d�R��3=�^�]�gekl��p^� �hGi���� E$}Y	X�$@$���EυQ�*�xl�`pjd��HK��Aq�:+oDd�r�qM�e-$2���:��ec����u��Q�{ٴx���,�+ܺ�qV}n�*����zU������|Z]������+T���k�O�BK8s�\)�Qw���^!���e��h�*����k����q�(D vz�큞���C��fF'��F�o��l�dCa[=�A��ޗL�]��]��0l�fS� Zhc��t�U%��F�� cb�{o�����X��s�٭�]7�F��L&M
Gq�}�N�x��06�ta�Qg��0�f�TQ=�[�%��Ltjn�)��p��o���z���}Jߪթ<�{0=,�2J�86�Q���4��p�&x[=����1�t�>\��b�c^g��2�`,V����A�/��i�,�4@�_**�tF͘���1O�#��k��C�|;�A���Ǧ'�Eh#`�Z(ʊ�j��g�V��fYE�-�������R�V+��[��¢��fj&G1��Jj"��qh���+���Y4�wQX�����Ɲ�42�O�V�iFN��;����h���|��H~���O+�{�cQu��u����	`6E
m����=m�p�y�=���>����q�}�ȑxN�峃ᘭ >�u^%�Ӟ��^`�ֽ��"��!4��I��F[�����"%����gXO����#�!Ɣ��fL�p��W_}5��?�~�* �^r<C�I&LX�e�' 
��&H�ۈ<��r,��Ֆ! Ǯ����9)T@�%�i#��-1|[:q'_Z�O��3����S4^�>X��]"c��G�ù�%,��?8����2 DH/���X��Z}�8x�`+@(����ʹW3�jY/
�ox��de*�:Fy�]�^2��,	XE�4U[��k[}V[��U�%V]��n8�<�����2�]���ܕc��1���W�
� ��3����P�'�X��3(Z�$����%��>��$QV�ƍ������d����l����S3TV��R)��H���Aa�^l��b**�M1�g�)p�����`�e��^�Bl75l^�f������fo�]طz�]����Xxϭ9� �u��6(2CXo�%$?�j9vN�Z �W���������԰]��7 (������h��N�;8��Q^Z���Upd(+�U"��.i�G��%������)[H�C<�'��`K����{}�!a٠l�,]H]�X����̲S]�qcоLp�I��4��l�������3� ���C`M�	z��=�S8�s�H?�9��B+�f�	��0 ���0��Zf�j����5&�tj�UB>;����y�����}0��=��8T�TP)4���������t��i�}����jP���*J�% E�q�մ~ga�ɑ���-nv�vA�+����v1H�7W�M����A��]��� &���� JC�9R���5�YX���wf�ؙ�	��k��L�I:VW�<@�j�������<��
Ǵ�y�TouSt�/����zm0�Ҧ���Z�l����ޣ����-��S�z�Б4V�G�n�����IR����������qa~�a�:a���]o�;�F��9���9�0v�a�����>
�M�%l�W�/�o��ÔZx:�p����i�z�q3�튕3 q�� ��s���D��y`��=�nܠ WF��_J]x3=J��q���DAk�� k�)3+�x���%��(�
Ə��n��|����C��JVJQw5�����Z��\d8؃�á����u��)҇-i��c�@o�?2���	\�h��'[�3�o�U�����휻�0a�'K��b��=��7�cb$3+E#���:��}NCH�4qE������Ŧ�^M�G1I��;�*c*Oz̴9� =V���U����e �
k�]��%|���"%LKV	e�m��l�F�ɟ��9elMXz>��y�=��j�6's��b�@%��-L��ء}y pP�|�J*�G+
��|�9������6���=���{&q~ş�Z cj+����d��n��h����=�Le�ձ�6�b�0`tQ$�˳XӔԬZ<uJ%����jm�����4M}���R}��@�8W-*�
vrh/������o��w�(t����������:4��>'�:HޒO���aqI3V̖��o[�$	��-.�]|��鄒
^�U<�N,��%&�2�U��ȭ[�$X�s��2L��d����0��rB��E�.�,��I���6wΥ���	��?`���Ҕ~���6�ô٘��Cږm�*��$����\V�Yjy�@�c;OX+����nZ[ҏ~�#�V���7{��W�f�a�xo�}"һ���˶�E55"�����!QC��n���`HbL�=����6Ӿl���}&���8�{��Y�����j�3���:�?��ͷ?����w��G���~�R2�FE�~�|�G�&a]�.T����C��i2�L7}��Rx���S��k��Xt?�����!�9�)�*��3Χ��{a<iӉE��Ǉ�3����5S䢞��L斁���a��O��'�+�o= �6&�5wa���q�Unj���+�A���� �tm��Uvh���t�Y�@O���guy���ۆ .����o�������h��5��~�v��\�����#侈h��j@s���c٩ޘĩ ����n �V���>A��~|�(�����}}ܿ������MMh���:kd=���o�o�ei��
 �� �3�JT"E8�������uF��``y����?P!,�C�ֶ�`� l� �l�l [7 N:��CI��X \��L܏������Y*ԿK�QD�@���2É���ͅ�c��h�[�����q�>�ީ�
bt�ϛ0�ZL��1���N�=�0dhN�x�¢�1�Ԅ���ٙYx�1s����ß�ͤP����T{���9]�W>��j����k��X.�׆a��pFsX�m�W���,�#���C����=�����c���N6Ѥ@���U�"�DKB�i�-�o<Ć��<٭Mm��&nǠg�ɒ�r��q��Sf��
��ʧN�wFs�/��fn��6����P�C*���C���Ū�������)Q�'�������3�EǛ3�'�_[5�5��U����o�
oVcc�������fM�ko�+mc�G�A��J6�@Ƭ8��l8R��ūGpb"?m�l����ʲG3 �%�H���B��놤�ɹ� #��3_-�=�`O#�s���� ŵ��[�0R*p6w�����A�s��~g�s]����D�����)��P�����wz��7[��o�/�jN�{�ÙY�`ɪl���Sv���LH������ӣ?P�h��d#��`څۅ��p���mSv'�n�|j�IGѝ��)����eg k����nǧFz�=�����hum�:��?�~����i��R`��B]wj�낎5f�x�@�3v���_��b��j��L��?Z}��G#t�:t���>�@����S6;���/���b�!�	`�k�_4F����g���#,,sheRa�m&��T�0���VطF�ƨ��{�fg���̊��鈡m�=F��J�b��Pi���=3��K�GP౽v�+�>��#9�����v����t�]U�Ѡ̈"�.�7�y_z�%곝����* �x�<�Vi?׮Ha�!�!�'{,,�������ճl�KƜ"��Z�>�uk��Pi��sڧ:8̶��C��|����}�Ű���V	~��n�̀x�y��u��@���݅�85��z�-X:<�mx��٩<G��
���s	ej����g����J�c~�>s,��K3@+,�x8�2��%x����O�I��1X�k�n�Y��4c�b��?��f���#.x��}����.�����<�2헆�����L��g�R�y�����P���_�S�VCh���_�n�ɳ8��%�P]%�z�o���������a�_��9��J���w��=7!�l�8���N�}�k ���EٟPIn�L�*z	�h\8��G�pp�Z,6k�G��/��R��5'�M��]O�Q��}�Թ;��ڍ�paȇ�����`py�~|����\u�l�%�c{�K�Z�$�FV��8?�F��EQI%�����؏�.ʘ ���y�a�ѥYZ%,j��*a`�*����ٔ�(^C�̢3������T��0"����ӶA�"r��K��Z�[
����e[%|k��I:a:�j)[�5�.�n���/�xmMB�qR��o�����h}�w_@�Q ȅP�&A��Q&[�|\0�0��<"ddRs�#��@�P��XöĈ�LJ�n3�p!�\��֘-��z�k��n�d�C�*t�s@�k��씌3�Q`5��Km#�Y}�U���������ُ(���w�~�ڇO�;A�,��N��Z �Ǘ��� �#\���1�����3��XD� X��1R�M����~���d�$��0U��-@<8�&sl��ꅆ�W�P���'�B�.���r�ZR̘XxMW�0�X7�4�	0]��8���y|=|4,�Q%���+xI�b[,�^�)��[���"<�w`�YG�FP ���)��gc:��>��؎�a&&r��K�>e���C�?1����ϒq�����.4d�$o�g���&}�8����N���C�b�%�Ͷ��dE]�A�"�Ns�Q���|#p���q�L�~�݅'���ߞG�%[��.�p���&�x��W��9����g|]Q�@��ه�� !�_G��y���3��|�c�a����'4�]��<�Y<uI/�B��Ѿ��@��# ����M3�ξ����Ь�i5MA��Whg��@M�+}�� �87~I.<��{�?� ������?'�`f�&l�6H�r�6��Et(�u�=v�X��Y?��k���)��:<7�[�0��i��903ֹ1�FpЩ3d�󙢂`�{2�ʖ-h+ߡ�Zq|��)�2�<�~��&�T�Nǀ!���&&pv�����Ȑ���f��|�&ߣǫc#��i�A��1�e��� V�%�?P90X]#��'��]]�1A�&l�,�@uN��o������UJ���F{�l�D�M�� N݌+u`�w�0�s͡LX+�I:��,�e�R�A9��~m6���P�b�����E[���h+��B�$����H�6��e�<W��u��e��iSmd۽��gIn�Q�S��yF^���%�0�)I(�ktF��s4z��������!Q�Za�Y ��g�)����X
2p��v����YRo�l���Y�v �L�V�i��`�L4��i*��2K�'=�'�n�K�2�P�ԴT�V�Y�{�,�aǵ�kpd�s�T�=�����Bd'�W^}= Cs�f���3�{Mj3� $�O�=J���dw9�<��k���˸�.�(�x���ga@ːݴ�:��}��f�1���^j��$k�˧?��,�z��WH&�i�<��)��9J1���*i���h�[���P	�5��,C�K~��H
�]��-]�7�jZf��6$��h/^��R�$PD��K�ǔy�	S���s��r����؍����E��U�O�N�#�qA~��'�{S� 0[/��Ϟ��A��3�0�l��d��	�T���W��v�G�c[	R�?�o�d����{h�=�O�!�h���*0+djPhG�����l�c\�(!X���2�<n㊻B6���)@�9B�g1-��3�9:t����x�n����Z �l�g��EGc�.�RG��~��y�ǜ"���ס([p���}�0�֡*N�>;���b�k�бX��e0VXA_x��j
 lM=��MC�����ȶc4(��I�����g%d̽�s�{_�~����dDF�ſl�
3Q�[�ȅ�%�	~�g���)�tٓ%4%�� ���<ct��4�}+Sz����@��d7z����3vꐝ>h�׾4���i��%#�޽�c����Bhg��j%߷���%�	���v�{����U{��t��4uRdjh��)`���3���.�v��p(�h�WuZք�܈�eE��\��vZ!7ͨ2Q%ȇ:놭�@��wI��]���F� ,����h�ڑF��lo�X�67�W�0A��mר�@-��Gj����d]A�=l�t��:;�nl2����nx�p&Wb�_���k!�P�}��_wJ�gG�Zt� jo��z ��#Ȕ�@���n���씄d�]����G������0�+V`f@�򌭹�d�p�̉�v����AFA� a&�3V�1��°;����pr�׵���5\�׈%oo�Q_顤j���kP�G��~��,���T{��y��;�!�l5��υbd�p&���u��Jw� �,��d��q���]Bc� �~D��]�tvWo�`�EX������ńB^y啄"v,��H��;+�aSQ��m��b�,����x��y���gӀ9�4���Rpͳr�8XfDi�� �PC%���؆�dY�[�"p\�3�RZ�:Sd��f ˜oa�c8O�MD���{$\����)���O*�����Q��B���D� n����VA����^�5�?7&1��a.�EM��χa�>/�Y���3D��}�O�;�[��2�g-�24炩���!�=������uy�A��	_��9,�Bʾ�(��*"W�[�����=ԴP� >��Q���mr�P�D�f:~G�\�4�+LP<���z/K����?_}����.�HYneh��	���q}�̌\"1!>��$S������iy]�G7)4{/�eCh� ��Ѿ����j��OW/Q���l̫�y���P�֮ ��Ej�ճO>��ζ�U?}�L5�� �M�+���h��P�J�'�F�ZL�|N��7I]�[����cܸ%K�~�cIxg$Ca�=�=%�Xï�K��L�/�H��{KR�Ƞ�֊����������;<Zf� �yʹ��0@l2���>l�g.��yzS���;/b�q�#e\[����t���O !�~?I+.��6��a���p�!5��N[����/�1��,5��W&�1OM�B5��ن������q��B��Z1��:�+����D�p��KĠ�����JS !f�0D����Ԡ�
�k�(Ay+�qM�J_f���ƿ���l�<�� �}�?�wr�`���;`��g H�O�0�9��^�ы��fh�z]�|E��`0��{���ʵ�(�������9�ڿ��ݳP�<�$�r�K�m�w����l�����7�g2p��1`�'?0�������'Xp>\}��?`�%�c:|;��t�z�}�jAoZ�;S~?�*l@ �Zt=�����@�E��#[I�ű����3�e�/"<&���H���S�?w��я�G�k)���/})�&���]ю�]�̅ Ʋ"^�2�du4������@[�W.k��}	g��|��atǥ��E�*���)t�d%�jR�]�>.Ԃ2KFX��2~<�%���˂L�òu�1������L\�y.���E���u`���T�A�~@���W�]K�w�ⰶ��E6�{1���3�X����-�`BP�"���)Ɣ+�a2�߹�*�L�fYs�P��e��]�`�i	��� Pֿۍ��;��c�8��j��"�u��R	,e�l+�Iϥ�2�;{� & �Cdq�|S������G�e�Ԉ�Eޱ�s�b�S�}����A?�0�:�����жm�L�0,ש'�������ij�y�.���抅4���R7O�/�z�����X���=N���i�{�+�r �"����|]����}\�v�,��*������^�&�/o�!�E��U�|.����T�y����T��Q���7Ihz	3�U��DC�p��=�I TH��̷"��zB�G*��"p��K4��P8x? ���I��X�"3s�͟��Ή�Yǋc��2pp�$�"�-+��nC��x��Gmʨ)��`�5�ű�S�Ò%.�
��-ٝZ���zb�y�UBHi���Y)>l~!���b ��E��I A�u���b�J�RAS	E�m�V��A'��,�|�D
l�N�W��zI�Ź���e������aӖ��>w���v,��.7�d����6��ѻ���(�*�--������2��X}Mx�Ƀ���i�%u��疸���:s��~��(�,�/�;�2X��r��{��و���� G�@�#�
k��)��Ufvmd�, <��u��4p�z핗R��A
��;�dfk�B�0X^��+�����2��a�8���n�(�s���V�;g}E�=�N*�gQE#ai���h4m"�B���8����aD�-��n�����L�O>IX��	�&�Ani����l�a�F��♢��Nm��R91��<��A����RΦ�Z[V&��AMq��{jfJf���K�N��2�wr6M7��
Cp�GP�^ȿ@;e?�0�B�
�MŶ�D��b�S�]�>#��oQ��P���&�i�}?��:"C�I���ڭ�&��s�]��>�j��J��,��48�lE_
n�{�2'޳����Gɶ��|��} ���wm�J�>��a+��E Ω7O���p�~tHGk�z�W^|���I�A����o�(T2.��2ӊ@����<�5�T�/�J T<��R��ݻ��B�2��d\�ä�1`H���;��c�3�t���F�����KN����L��0��2.����`�V�z�f��4���>ct�,��3������b�q:��RȄҷ&�.@ �iK����1SL�L&��+:�����nX�66�Y�&l�X~��*�"����{%���aC}�8��@[5B��v��,{�
�� �f�0<|�ӹA���Q뷢ߒl_�@u�%b��M�q���^�6����zX;N=&���I�L?*6�z}9J�" ��2t��˧��B>[u�2�:DKy�Ο����gG�'O�}���C%����7i��_u��@��B���ɖ�:��\�!�Ġd�)����Y-w ��0�u���� ��"N�j�� no���yЧ��.[!����wz�駷�O��?r;Rᜠ����
������N��k2��7��8m[�9�^xQ
":ae�ʭ8��	wt"��ޚ���Ը�;8 :|�b��Ȏ��)��It��?�2Oz�5v���´�T���ɵ��<�z�]�ev���@��M���S$�)���wւ�YX�La������T�'2�����oR��Zک�u������N��@b~�ڃ�L? ���0�2���ϒ����U���da�x�8�r5��26�*���Ta�M\�mP#���h�����8a�yw�?����5Hԭ�E��/��ޕ��/���	�����30?.v�Y�sl~I�V$?�g�m��fx��u��e!�X��]tZ|��5�]5:�l��s޷ H���(A�y�
���C�%�8IקL�A�Wĥ|�s�,&+k���L5@���`;Uք���K!�AR�:���yt����
!ڟ��'K2g��.�zC/5�~�Tu���}��9fܲ��';��]�2�� �Q�v����<�|��X��qf[x���$~���V(!L��(J��e:���D��;_�j�)?}�8\�y��B�t�N�"�U!n¹��z�N])J���u�������$��������:`6e�̾8�6]%m:�d�{�O)F?��9Z�#���'��Y��_�����J�5�7D
�Z����M)��Yl��%0��t]��9�ŐU2��`?a(>165��Z�ܯ�燉+q�~�S�,��� y��� +nj���&!3�=
�v�>�����H��<^]��FAyP~�_!F��n����b7�Vf���NVvgWa�l��2 �l,�$ud	o
�xOk����I��`:���&P\��P�@�:�`fp���R6sP��:a&�SZ����sc�톙�����g���6Џ����Gx�ށ����:׺(�ocÂ�z{�|�����2A  �wz�7Z��ҹ-��-�S�(mxL�OvL4,�)��p�zF�0)�QpPeQ 9I�0�+@(��L\%�[�4U�5��݄faNNn����%��ָ�u�e�<{�,`ٹ�@�g�S��?��Tt���q���d�.
P>���d=�����x��;��u 0���e)���;��~��̂�X0#;�a��]��P�z?�OWϿ�<�u����K��1v��b�x�e�FS�e=��f���ٻ���ף=`sgo�)ٗ_~���}���GsmM����������'��~��e�tBNaLv�Kߴv��.����#�gd��%���{�I�ǐ�疙�N�΀�"W I>]˘��{���e��4�;���Ùܯ��q����s���=��d�Al�I'\3�m���&��/���]���Gq
7Ķ�j4L�,���L�w�
H����R<3��}ֹ1}3���1\���4�[�Q2�̮:G����G�.�VWp{�uz�tt��Ƕ��"�w�}����=dp�#�v c��7^{%��f�q��^�*x�:�g�;�{������-� ���d~�>�D�UC0��#��Vg��0�Sm�Lm	IglY:A�U@���X?&�����C�t����>[������_V�� ��3O֕Q��+���M��~��R�k�� �Q/���!z��AJ�/���5EYe����@�M���iҥ-�0SX��;Ƣ�V��K�Y��F*����r,���&��rnJ��v�X�F���S��}:����ù5�ܶ�:�x�P�,������M9���>Y$� !� 
2/�#ZU^�����x �}$�;D-<2��O�+6c����8����e�4tD��`sի�RD�)��>x~= �>�>,Qa櫦�L�]��%/����v���F�-��l�9���\�kl�vP�R����U�ϕ�	s��Z�i[�@��2)b&��AA�m�����dxV4���M@D������������n�a�z�������r5}_9��Zp�[���3�}G��������ڊ�,Nm�ĺ�M��Kg�T���e�A�Lg܌ر��6Mer&�v�Q��"�S�V�GpL��"��d�4���,�����Y�o+L�g���,@v����H�qa}��8�³f�T)"fpά"p���$���LH���=ro�$YG/��v���on:���O���׿V]��0���ԝE�B�j�ԏ�#�c��t� H�Xo$+v�O�d���z
��AĲ����%�,zy�j���P{��Q�Ek|�h�&X4�=~�^v�)P:��hQ���~�_�w�| qOu��43��M����-��|1a � ��rӼ��t1���q�gAT��B�w'��z�x��h.�G�M��b~��U��O�V�1ɏ`{�bz�n��>XR����I��C�vb�e{��4��#���%�t��%b|�4� �c{��=[�.�]�`���Z�w���0�d��W��ϳ&c�v��0[7��p��\=�0ڧ9R�YTJI���P[`Q�N��ajy�!4�����NW��%����f:���u�^',|��t�������y�z����gj�d 2@Ϳb�Z��qJ��V)R��8��9׀�T5�#I���?_��_��`T�0���\�fa5x��Rp����YP�k��������l�,u�gMg��s��3;�u]�x�� ��7~���������Ļ�jO�V	��g��Qlx�L�e��`���k-�.��h�6�'����\[ �ʂ:˴���;I��-�t,�kf�20���8�[[��Ȩ�~�,@���0t3�eEjV�zYA5a%�p����bWtuE�����1aB��� �]� *�5����d�	}�-Vck�y��D�bAѷB�<�9)5���t�4�b���p������0V̔�����_�lUGw]���r}&l�^��2�jE��P��˼���2�|!�Lrϳ7muxL�]&���(b��GK�P����)�6<6׾��}�����e��m� ��*m���8}'�=��YF����e���b1�(�ͳ̉��D��.9�(%��fZ���綦(7 #޵�9��Ru}wp?���c0B�h��WQB���m���	�s�Q (X~k�G�Pov��?���:�,;�)�� ϒ��sv/�\�Sc<�]�u�Qs�6��7�Pݝ�SQ��TZ��βN �
���8�
\�-�1nD4m�u?P�NVZ��9Dq�Ʈ���)��Ή�����1ˑ��	7����;'�`k����xX9�J}K�����)�3�n��Z�n<d� *��VX�%v���K5/���=P}������_(^7�fa�&�x�r�J1C�KM
>	���+(q"�"��d�̒Jo��{	��#0���~;�^P���nf���	\�S4����<�t�qa6|�g�쵒ʹF�q%���ǐa��\���L:Y��g/ׂmS�K��%d�k��ȲJVd�\h�3���'lv��9��R��!Sֈ��k��X̋g��d�ɘX-��5�� ��zoև��1�EެW�
��z�$��PX]ʺ�Ո�@b	T?���?o ��S�����_��>�n����i_��ɶ���vFl��N�{2c�6�sj���ʽjR�k7�`	��?��#�'�L�e� a�YZ_�ۄ^5q,���QYa,��c9H��Yc�{�'�~�:y�$�Z��n���?�Iu��3*K�dCf��fr}��Bʋ�a���$�=?�1�11�����l��q���[t����z�dx�T��o&�obW����0����mA5����|�+l��f��?��k�o4��E~�x�_ k��э���)n,#m������٠,����>��Gi������`���%0,�.�p�~ ��2~8���w	}z=!SjM$�Q��g&H�ڪ��B@��+�jAP�q�V���6y���(c�z0yO�A���j�n# �Vئ=7@I�*7@��1���I&�����}�MeG4U���q�_`��ƹ�N�!W9��)�3Lu�V�hB�0g�8q��ͯ�r�V�0Fs
�}p%{-�;��[18q'��!���A�ltt�NXˑȠ�Ǩ-{!?��}s�E��N���`�QÄd�=3�n� �^�M3!���a��c�݃s�����/��	�x�*Sc�y�8��ڬ�y����"��T̴�$jB;��טɫ�P7g��.�WG�ab�&����S�Ō���SO=���d
D:��Ҹ۱��������,�:,�n�0[�}�]��.��5�5�f�w��e�`'���C�ӵkT3H�U� !�����L*ڝ�Mj���kdH�X���$�;���ŔRx��)��x�ÊP�$�4�K��^10[���^4
`����1TքH\h�%�y]�un6�� ���� �a��{dgݤ k/��N$/�9Cm0)4�f*����@q�����*��N��Jޢn��7��y�>�>��\0��,�ѷa�`��X�E�#%ؐM�
6�F�Y&`q���^�`N '�3�ݶ��o/���}]��L�{<��/���o��)τ2e�h��<�n�i�@E!�L�e�7 uuz�Ԍ��M ����|���#|{"�@�sj����]u������p��4g����筳�Q��]��.�	-8�+���Ha��������6Rv�������G?�I@�!�UUP��^R-��������W:vW}�c�{�u}܏u��M0^�9_��0I����������F`���jx�qO?U�P�s�7���s��r��a��b�Bbz��!7�W��d�%�L�(���l�]B�%��?�:=d�^s�e8����t�<��	�e��W	�� ��]|!�r<{�����ćYX���U.��ƒ1��]AC�3LM9�%�����;�vt��#n�$�Fː�f�	�҆�Ϻb"	��l4�v��ZДOn�I#O���uo�q�ZF�?�2]� q�n>�0ˡV �I�)L��ة%���c��\��.c9O�>�>[����_�l�.c�����r�T�� ��{q�vc-��������(��o�W�����%��G�F��2�9�x0�?�J���!�tbs��׃��0��Y�ɒ¹�6�3]�A�.��dJ�|t@ř�	ɝ��{�16��D��"���-��n��dV�Z�S%Ka�{�,n2EI�E�����&fe�o��C�~�[�bbZ�>B���;����,6ㄉ�~�b1��e.����j��;9ʈ�%X2M\�������7�[�cj���T�Q�¹��o�k��=_B��,��H_��u3��W������	�S���'�N�jJ��2�j���b!w�7<'%o���D��0�̝��d�P �fA��ͱm��(����6Uy�t~��ӧO�M��}�(�t�s����q"�z	Fi�e��O޶w��mCqܖ�������� 6�1A �,�`�s	�4$�%��cy�8Uô�������|�9�Y���Z���^<-&i�t��hliiA�@I��6`T��������q�o%��/�1N��n��e�FY:���;�{R���?}��w��jt�N�3<g���,%�p>k�K�2j�n�Ȋ�=��hKC��4iV�N��M�_���ݤ$��6��0�2�H��/�z�����їd̻!���`F����%:�Ҋ.�����#$짌�ۀ�	D��h�a]�	r��eBdi\{{<��م��x�%nBL��#�������?	���ۦ~�hP�#K3�X�MP�
|�U<.*��1̳���k��S��'h�� 	�[�|+%ڋ�KFSsʋ�6t��`�l�ٗ��>�mu-x���`
��`�
PP|���R5]��V��N��8A���� �1n�i�17,er�
`c���ݦ悡O�Ir3u>f�m3on����ғ��j�H�}�xz��ё=8����� }�� ��A��٪��dޭ:i�^
���������~f��>�!\�3G��:�� �	�Q�M��@X�h���J�;�іv�Z�A��;�w*Səf)0!�M���L,�	ۆx^8�m2����n��6";���ٮ�vU��T{�{Ȓ&�`r�Wg�v�O_ұ�� ��q���;�5��,	�?DQ�"LƮ?������j
�hV�'�?�)�Z�-{��1M�~���Jk�!bT�8�X���d1�����^�b-�)��>X�����iC%�\����;��e�r���Ņ����@�s�"m����?�XB:��	��E�����s���P�3�sѝ&�����<���,��kr�gJ�d7��;�����Kн�	�J/"CG��|�0�,�,�@R͒����p����	R�/�b`��˝�*A!�K�2B /?S�;��BV�ЗL��l�k����^/��t2 #���|�k����{��aS����{���2;w�*��z �;e1U~'K�g�1�P7�-е>���D��w,��(}���f��g�.�^Sl�����'},�{�c�KpV�82������"2�P��4�� p?�e���}L}�@D��\r��-C#�Pw����1I�K=�R[�~)��5�0Aq����~ ���k/T���ǪO}�1h��w����E�!%ƹ��(�5][���N�z����|vW?�ُ)�z=�6(<K�H'�@ޱ�N�a,���5d��YH +��w��!�"6a�b,ꗓ�C~l�¢���Z3�\���ky1t@���fI��L��c�X����eY��y��1���TG��q��Q�a�㋰}���pˈ|MQ[�q�%�������X�-H\��ý�V/[�]�l� 9���k`�mH����#R�G����xeѭ9F|[6l{U�pY!Y/7���lv{a����ۥ��(����G�m�Յ����k�	3kIǳ������a�$ [�1����aB�d��'{�ﰅ�5�yk�ݶ�Lْ���<� ��>c���Z�6�L�;g�;�|pwǁ wkd�l!�m]"����±Ae�������>p:�Z��2`��nb�G��U:x����~���",0R��u$�/�э]�e���b�U���L����M�ĉ��~�z$*2�fRAWt�m�j��%b^\w�ܖ�P7�߆ԪU�Xf�4�N�Fg�m�ߕ���g��u�����{�@����� j��Cg�^I{�r|��D�f1H{I�1�b�D�"_�]wg�|�ɪ2u�Іl�� y�6�E��,�����q�֘o&��$>���¼��^{���]BI���x�L���Y(z������I��+�[�����;�;�*���
 ��M���l#��P^��s�*Z!˧Q���Y�2�1L�,CwO0C$��6KC�]�0�KS)
9FJŦ������}�א�?�N�-�������	 �)3����n�
�����?�O��=�`y.	����ګV�7�m���\�`����%���C ȳ�U�)�a��ٹ�w�4.�lwU�x�|��V�X�O��<�6=JL&	��Yߐ�պ e�fF�.�L���	�j:�{O܏�l���1f�=_���[������Ƴ�����&g(|J�f\*��d�D���p��Kl��"����?V#�=r�q��[:���r����Wł+��k�_c�W��q���$��F����D�u�h��3I���"�Ï��v�4���R�h�<n���Y�����(`2�̱c�i�1qy�(l�(�1`h�1�]�% �>��A�������f�ᾦR�O�N�9������U@^R�-΁)��G��Y\zF)���������3׬���N������A~�	(ʼ�=p/���W0�2�����}��q�]��	w�7P=tx����������߉H;!��پ�&���׎��Y�i���E�(cy=]�:6�$B��v�dMX�m�.s�E.��m�5jW�5�!�봎� �	��ƀ;� ��Aw:u�l�_��������<���eV�a@��6�9lm�(�����em���GvT�8��믎���b�k�^���Tw��,8w@���3r-�h��m'\�me�N'-���,�h�Sg/�	��իG١����Zb�o�V�oN��'t�Ԕ�����R����o��T�2i�{��S]�~�pDw���τ�y��/dg��|fb����P����V�i��1����e�8#�s����xY5C1s3�t�ч��>�фL~�_�z�	ءW��+�~��L���ɘ��z6un~���R���!l�q�uq�j���<a
ɲc>C(�̖%JdQ�Pg�f#���7~EN�����Ӱ5�ag&�����'���	2�L?w����Q��=�) ܏�D�ư�)熢���/�3L��.PsɇN<T�D�5K�䡇�v�
�����/�	��T��L��,���:R�'tP6������������?+���H�pU��"��f����m,X5\�9t_~�G��7^{�z��i�̞�Q��0�뱼�=�9�;����.kt�z��7o	��(8~���O�)w�GA��L��c�?!�8�,��?��hziC�#��dS�m�]��Cܫ�y;�\�E`VZ;}��n�������;�V����Y���x�����������_}�o�5M�0�	U��wc�A��WJfX�>���4��mt�s���9��Y�AP��u����IHT7� �������`�n���̋��03	�v)�L	�Ol���iBOk��`>��}�E3檀F/h�x��JP�1�1����r=���Qt!��R#3��D|©��q�0P���8קV�4|ƞ@^��:koay��?�9�Z�pu{�C1�d��gm�eBA�P�\���J�.uW<� =v��_���!Q�c&�tb}Ǥ�ӨD��uR�T� CU�c$����g;�3�u�����{��gu����=�V;� �=���<J�[��̇e��L��߲T�Mj��̐�8��:@�c��#@�����pk��c���6)��deoz9�㨽#x�*I������(Ă�Nɋ��驭�UbFR�G��Z��� �9��4�����v�z|`�z�h(<I=�{��w�~&8��B�a���wم�����-��Rs��己sP����V�6�:��Bp��C����������Yv"��q(�;��\5�,����bnv�j��LB�hW�!�]��w�Yu
����0	�����+\�!��C�ؔŶ�)pk�\��W̺�����.���eMQNlfI�j���ZN��� Ν�}�e'"%`e���'� ���%�+��(bA���q-�)�:~�\�<B��_�,���f�-=�/�ĥШ���~F�A�)>���6|#K�HՊ�2WaEԩ�}���
�b5
�T���!����rw:�;p��\�\ ̖��f`5�FuAޗ�I��\�B��¹G�Y��̘nԂK�r�m�*@ݓ`T�Fo!w���:�5��(\��qO�q��������_��5=s�t2�y��&�r��Yc�Ȍ?��,[^�+��E�PV623#]��q2�]\�<������o�q�[Hm�a�% ���=���3K��H)��D���1�s�b�H�?���C�j�>L��!�����y�֓O?U}�S��.�-T�����BȴU�dc{)v:��Dh���"���1׬S���/�3�F��Ym�� �`L6Ml�~��]�����PM����j�s�z��w�uλ�oDR�G}�Q�2�Ld�eI4X+p�d^ؚK��LY��)@J(�v��^͘��ĐS�AP������D��41kTۉb��FF@�>G��]��3�ŅY�FjV�$�|Y�7CE<?}����4]g��.���4���f!��+ݩ;I}�ϸ���:��qiJ��Im����0^�67r����G��L�Ђ:�+�WH�����V޻�z�pou/eP1_�"l�:^~���W�Xt\Z$~X��҈EP�秮���Xt��aY:H�Tc7�	��Bw,s�~2���K���k��5���o�Lv!�G��NڪO��Y��:۶[��}}-pG� G<1�)�8��[����"Ƌ�A`+���[���;��Pr�Ȯ�C�[�܀����8t�(���R�gqgäh��	����������ue��tS�&]�� ��6+<3�֥�	'9Z�3�M�l�,0�\�D7�Ĳ�OG����_�3��c�����F9��4�^؂g>�\�M��U?�r�o��oe3}��Ǻ?��ܧ�����3D9�&|�І�2N
{a���O=ɢ���\͚)��cOj�P%��;�V�r���δhC6==}sScJ���;In�,�O�<�(�ڒ%1h{�}tUG�r!7�3�P�P�:ʲ����R���h��ЖY0���`d/��g�c&��kA���J��D�h���G��E\ք�bT�w>��.�N������3��B%0��yv��� ǌ�," �z�>ϢU��,�O���e���m�נLggK���n���B�j��G��!K�/pQ+% b�P������qǛ���� ���e��2~,�����㣏=V}���5� df�e3V���lmw��F]�ѽ�>��.�-���%�H���"�ꬱ����K ċd)�(���_��}�����'�e��?�fu��2%�Mv�J�`[��%+o�S�6�"�� � ���T�%�W	�
	/n0���CI#���ă	����soVn�����27��1,��-����+�@�������a���!ľ����V����q���6��
ҷ� �gA�Z��b��<�nX1!�M�cju:�w�A+�J�����s|斚u�y��tcԅQ��7Hz�*=�����ff�L�Is��5BZ��I�E�����>W.�iE��ٮ�yfᚥ�=�h"���v<L&+��E?��dXHo��9#��M�D�?0h�������j�����9������_Oz���ڌ�h�DC�����/p���|9����}$ttP��²���d�mT��򴫙]�%ꇭ��vY�}{#Ra�%q���j�x2i�}}-pG�  қ�Vb�����A�
���{ �� �а��ƃ�ՉC���������o��CP�n2�dW� w�$�At|�es"�lj��X��Xspu���Ę�An�8�f�%�C�A���qp7�u�e�QD�Z+�	=�Z�Vw����i+�t׼
P�e�84�=\]�x%N��<�\�E��^}�z��g�!x��q�!�WzMyƥuΒ5>JL\a �x6�L���,1���zi#}[L�]g�I
6��IJx�%s�]�}��Y��l�a�����9X-���J��lL�ZHs�VmWXn�'���D�2"���6�Y��e��4��D� F��y��aؐ�H�]K���ژz�	�ș�%c��gf�qsj"`� �|�AOYDٍi���z��8f��4d)f�e�d�}�ݴ�%'|ӫ;`�\D���Rc��~f�Y�M�*��3�5���c�)�,�Iᗮ��d���# �Zo��cF��3�wS��������m��y�CS#��D0�$BR2��k@�,\�&=�!�"�7��_N²@꺾�qPq�U2���z`Ĵh[��{_%�d��~����}Y����E ���H�7T"�T輇�5L�y兗���x�z V��}g���O^��`�j�� bi��d����Ѫ�6�g����W�,�v=� �G�0YG� �g�A�3EF>�TZ��W' 	dM����B�yɮ~��ӟ���،�1~Г���|��E�aQ �7̥������&��jS^	�D2{1��:�,ӆkͩh>P{O�]�Z��%(�!��F/8�����Em
��hSù^�������1y$��8M���=i�+��!l�>'��<k�b�q��;)�L���|9�����{�=1����-" t\��`�cm�,���|��(�%��7�)�z|�^IS3�Y ���g�]k��'J?�'�h�
�o3ʺ�:Ԅ���,�B߼���|�r$��x?�v�1�|���f1�SY[��I�"6��a���wk�} (}�:��?�f����ZI+2B�a����.������y�����g_u��(z�>��N�06�B�rr0ׇrgK4��Z�r��2�S(�2Q��1��Np~�Tdoe m���'3���$�8]\&�us��~ɉ��1w�e\|OՐ-v}�tm*`���={����>^}�ُ�k�A4�fu������I!C�k�U���j'k��+��C�������8f�R�]��-��,�2,��"v�|?`�>0�<�p5M��g��$���w�@X��	4#��c��+?��0�/�2Ȋ��4
�s�G�`�y0��6�F'b1ɫ�Ԥ�_~�������fo.�2(2[��?L�v����E�����U���>ׅR_�?���.�� �T�6��@F���H*J����m�$S�!	��,�f�dٍEhw�
�5��%3�H g�0Mq,�(��@�E�*!4�+���7�!��<�M�f�јAr�}���۝��j21�r~~��D��EM�6�ax45�l]�ڶq�n�uP�W�>�h�6^�!1��fj�M����̐�ٓ������5{'�_��Zq�#C��%�xps��x>�ߣ.�����T_�ʗ�O|���9����_~��t}�Z�v[OȘ7�;�{X�P��<�-G��,��6Q��L8��[�]����˼Q͘Z��=w��$Y�	tћ��;�8i����Bٌbŭ��V�����F�d59A����z~vN��p������j�U��ϲ��4��'�4nR�[��\�wg���w�⦫,ڦ����v�2�^M)�8������dL��~�️|����$3�i���.r��@��6!��-EWĿ�hSCJ��M_k_��lz`�/�A�bC�B�!�E���}'f���4���J]�-�[������N�8З�� eL��N,� ;u#�>i���6�1�g�Z�8��vJ֩��tq��"`M�A�D_ue�2Y�0B
�YO���NV���؎�L�Um	�w'���m����w�d�cB���W�a�}7�5选\���B8��9V=yϞ��ž}�RH�A�a(�2Qgp�4�wzi̚��3-�M���1��&6�8�b��s��W�C����chzڔv�uN�~�)4[A�'\y�͝���x�;p���գ�_���\=����~P���ߙ��0�LT���Aq���bv���n�/�J��-�}'S\�m�4�����1��~JFX�U-P?Bd�~L?��/$�L��Y��#���}�K��Q��"q/ ���lH�c9�`K�~8V�����&"Ő����y-�yD���_S(��%�aڹ�TM���D� @.r= �n�}����hY�I�9$m����,n� �� 3���Him��z�����������=
}`��7�M؎l�Iz�W'�ED�����%��f����^��u��SEЮ~���m�ˬ=�T	_qΣ�������Yl�h4.ѮS2Ox#Ϻ,jsRk���)�<�+}�=�B���g�5�Ţ���IX�@�a��}�z�X��fL;�lbi������a�Z0���%���� ���W~����_}�;�!�5v����.v'x��V��'I�X����S0;�(��%,�L�����΂n��F�Y�Da[0��Cq\���P�Z���	��kv
_������le��,���fd�nѧ:x�f�Y5|0�c��U���e0Kvr��Ȳ��R$�)-cY�QC��s�B�d�(���)#t���O�D6'4� ��[�.��D����V�}d�Hdz�O��p�� ��DaV;���碌z;a��e]��l	�a7�^A���8��㐑��M�_�بl�Bo3�uҦ�.�9=������Cp�^W�:G�آݵB)	��f��C��k`L-PӮ�қ�=���.��x�PY~����)��H��X�YѰ]�d[�x�� �`�,����a�j����z��������d��A:�3�7eNB1��K�/�I]�7�S�h�t�QR*�Wm��al��������1��4͓k,�o�����1v~�6���ܽ*ioń��C�pa\�[ݘ�A�]+!�������p��!6?����8U}�ED��?�)�O��ju�}���Z�!����,���|_6!Z����v1jgn��w��DD�B�O�,ګ,62�<i%�*�~V";�&��\�~5{?u�dT��j�F���v�;���u^�|5�z?��`��y���d��>k�O� {aU��i񾬌~����2g��X��/yݳeJ���3W�����dh� ݠ2�"��w	�1�{���n �`��	x?ٮ��e���݉(:SVwG��}��=�(��%�����`�N[��	��Ә.��ds��a�y�^g��r=f���-�mÚ)n�*��j�鱺c�� �� ��y���?w��6tx��P��2z��y�K�م��L�S���0b3���rmӯֵ�vB�㽝=s. h��;��웯�F��P��/}�:@������B��3Ăn�/eiL}7.�Av����IBK<�VC%.~.Δ:0�=��q�udŪ4lG��J_��������DHI��zSђo�m�H넶�I�6�D��s�
��qT%�=G7b��|�d}�	�t"���^��z����)�V&!�#ty�;O�f���>���f�P�Ly1��V#�F�oP0܇�����-�����8�b�5�`�S�M����2	���nB��*��1`.�>�`�Iߧ%~���<V �`�[�&�4s�KT�d�;�	Ɇ=)a%�`���Cdݳ�pb?��h�e��#�(Z��[ l~�f�;��u�3�H-M�g7�Y�� ���{w�ڦ��4`{�:�{�6:;��
�C���yk��c1�p��������1��f���r��e��VE4����!v�^*��T�ʮ���N���Ix����r]�L;�M>/ �ݩ��' *[�2Q��e�Ɵ�ְa�s�j��H�]Xq�fݙ�{k,��*'
+�r����[#{a��~�����3�ȇ����ߤ�����!SӇ1�����W����;f|n8��"�
'S�4��>]�~�aя��3��S�タ0���)��a2\4	y��\gl��:�[,L��c�^��Wa���u��R0D�t���4]{�:�A�*���a���u7:�7Iw���uǶ�{S��;���nJIo�,w��@O�	� ` �<e/`�vY��k�x�bjo�SHv
p&p0�%�x�I�F�K�SYu��-e���/���$���F;*��6ם���Rv��|o#"�����g� �ŉO�W���W��V�1��w"�����d�|��ܓק��8׼��H��	���)іn�!�˄8r�fNeW��b��^�|�JIZ��k_�Zu�=0j_��oW��G����[��^u}bN1:��&��޹�2,�N�5!�0I��!�k1le�B[����&�S+m�YY��K�*z���>�=�(q�f-y?� �&s�^��s=�ס(�s�F�LxN�c�><��f85^:ދa4�V�@X�땹�j��y�6>i�-Μ�3VߢF��XjV6-�`H����nLҟ-T
��9�Q��2V]�7 �[x�l���L@�i�u�4�܆^[b<�
�k��
�Wh�Fa���W�Uî>0	57Ujqj��т2mZa�V̚��:��;8
 ���'��	�
d)����-P�~o��޴�i�F*5Sd�({�&�̇Q,��C��<o0���&ё��6�up� �)S��3!,�T�l
�>����)h�;
�=ɐ�.�֌�������u��6����H��Sd�޽�������	c�ݧ3����4=��${L�o��e��Ъy� �"�s����ꙁf�H�!h�����Ut*,�Z���=����vJ�8ƪ~#L��|wj���`ܸF��Ǫ_�үW?��I5��ZUX���NB[�._�NG}��u	��@��2�a� J3��膬����Z��� +T�_v��3���aFR����Ka�d�|�b�,�a�,� ���43��9�$�"�c�w�L�2@�]���]��౽�E�`y�d�F����S��ط�E�s_?�ɏ3�j���5�$���
.��~����FM{��Y�cA������u@V��o�A��+��p���.@�B~,�@�K�n������>qc�����p� %&�i��U��|n2.�����bC����ڎ��U��j/<���V�G�M�k����}���1����O��z���҄2���2�Yk�����ɒ�h@h�²֕�}.�	S���v���M7�Lx��g�%v��{�~��깧��>���Qz���Ͼ���O�����!1n�d`��J�tw�t�K��~%�g���q �7�La���#� G�cASh�Ҿ0�۵�ڼ��[�ݬ�%�(w�p!�Y�Z|9�Y��������#�$87�'tC��_�*:$� TI�O;5.���9)� �� �=���D�'�S/޲'��.��;N�����v�-�U"��F�k	����,jt�g2H��e�I;���Bhp]� J�
@����d�c^�����G�Y h���sѢ��h�M5A:O� 2���x~��c#`�7�&nt�y��1�l�`{�"�ɿ����+��gb��o�7,.#��_6����i�[�дY����XDQ��
�E�0��[�τ�u4Xޘ�}f�z�0N![�J���Qmk�:�m�j��z�[��A��=���?��]����D�Ů����cG�� ����������O��1m�W�	�I�]: ASqn�S�l3)�������^%	s|w�eBsg�a�Hu�����\Fٙ��jM��t;:ـ>�#22�@��L��x�b���\�v�B�����W����s����%h��,\+��Ъ��d���7��1m��֎ ��ֆs��qW�=��z�TO�{�(�w�ɹ��ڇ̾{䱤��wߵ��eG&3	.jpȽ�2TfI
�u]�u~& U�Rm��)��NӴ|S�,��KP%+qp����C&���0R�}����c�fGfH�`݉���#�6d�ӟ�,:��i�IU�?���f0u_]S�=��j*�@D�C�%��K58H�H�1,l����i?�S/����Ȃ�M���l@1أ_)@�?O�<�~S���� �k��]c�H6sL�r�t�݋Yh
���M*���k�\>Iy�����l]|{~�kWk��K��ktz�> �]��R�gj��݃�����˿��b�����?��Ä ���_T?��(�U��O�`qN7;dP�	)-p�,^�V�$X�� ^��h}��&�(���PL-at+��VBT������E1�����=U�!�d&y�{`8�*�5�=c�6��&�z�l4��-�f	x��F�{&E�^I�hD�^�`(Gu�|@����o*k�8����&kέ,D�)�7D�eΓ�歺AHΑ!j��q�aZ��	��l�X4�}��=}RJ~��p�ҝ�p�!:����ׂ�+ت ����HM����axV�r�A�f�{O�!60�ZΕ&od�T3e5���D ����?���v��R��<����w�{��J{������e|�z�i �����UV�z�!|�Hw�o�0��|�e�>�9�bI���@Z��A�zz�h� tVi_���g-�|CLh{a1�b���G���3,�L�0>�,j���2	*������;�|7�f.)���^�fq�������{8��q���U?�qX�v�������x���:?��v��+T�^��]������!:�AL�N�E��_�����SOQ�j&8CR�]LBn���X�����>1
�p�U�"����dP@�s�:�jC�����lB�G(�a�E~k�݀0U�Е�ȅX�CO�	��<N)6
���K`$`L�� �c�E�c�o�C���L&G�e1�!�'�_ i��;MA�I�d��ߑ-�G�m�I� �p�٬XA�`JVF��+Ȑ-,5�*w�ay��(l��E1�L��G��V]��<p�bؘ�jo ��=�b�hxl'�
FEq�di����V�k�YB���0��W�P�Ah�о�Q���f�0D�uG���/0_�;>��CH��2".h�Xp5�%�ٵM�΀�m|��S�*���kaA5�S��y�K�E�ޞ�Ї��:E�㷿���g/VчlȰ��ߊ~MP`�f,)�e<�`���`% A�2�^�jX�,�Q�#�W�\�"��W�?�å�0��a��\0�#�)��y3F��W䵔���a�H�P����3c��H��*�%50	�x+E �,�){��z��bj��&J��մf+��X3j����3Ml�1����EB��$�$k��,�:�֦����؆֫���K����	�,��nx-MH2� ��J��v��[q�:$3Һa���[�$ӊF]2>ܫ 9@ƿ,�o��(���
�(�nf���0Y�y�D�_�ne����g�sn6��}�;AR��A �g�q���~�m��E֎[=��`$�bf�P$>�A�������,�ٸڎ�-�0�L�w_D�Q ���I��2ѢI#o+NuH���dk�{W��*���t�N��,��ZQx�$=�J�Vvv>���P	��"-���g9S��L&Gf��10�%!2�2���G��<��.�*��;\�)���hA &b���0�'c��������Dtx�µ������?��ꉇ ��]����՛ܹ+���+_��8���?����!�h�����YE��Jcv�}wc.�u�*4Nī0f�
��I݌�i�LlԎ�fX`�x��,��,ކyl�drqA�N��,��uv�.���f�j�Ƶ�[6�!�P���eh����ˇ�jZ�~P�#dO)?H�(=Ff�3�((�p��S�ݚM�9����4����f�޿܀e%��F3�ܕ�2��{X�h�]Cc^W
���E�k8w��/.G#c�K��w�a� ��N?�E��7XUwQ;4v�A���w��2@��@Y(�糑���n0o��:�2%_�5���Q�I-���]à
��.&1�D��F,�(S�so�����f+��h����S��7~�������:uẕ������uA���:"MX�RY��Q��V�e���]Ͱ Y�^ U
��������,�k�&n��,�S�Lɷ*�ɸu���
�y$d��?�sY�	s��Tp���I�Z�ig��;�2�%-��"�ĭN͓q�O%��c�V�M�O	/L��*�q��)Vo��������.�$`�,H���HQ�1v <���8ڢ.���Y§)4�,R�	[���ƙ���2E�}��vMن)`mg��^��yB;�g��f�i&ia�8hh4���v�G���ܣESk�rAf6m%�߄aӘ��z�e�nKj�(���=����-�Wҽ�yi�}ci���y ��~�op��<.�&_���}݆�d_��N�I���JQ������(�n�"�l��� �I�L��gsd�0���0<��:Qab
��_�J�^b(���������ba8�i�Q�|��AR��ؑ�PS�e<�����?��&�X�D��F�Qb��`r&1hK�s&�v�w���b�@��]I�|,�����2KƎ�UvR�F�W/�y�t������k���������OZ����uj3J�KWQh?�6L�Vp���D@!�YhL�R�m��`!��.};Y��;i9o[�ÅԌ��1b�e�����.���/�G�����~ng��7�����@HF���0�n=��q�� Y�"�
����֝��xW0������DR�����(x&fՙ�URͭ����	���n�P����,�0C:�'��|f��#Ȑ�I1�YGF̾2av[ �EVa����w� %}�R�L!wa�6�\����YҋYt�~k�]6�,H����\�L�6�c����~�W��9�6g7׹\���O�Y�>cş�X�ؽ���"P���kZƀ��p��Ds�yB�B;ڮ�M�����y�r6�u�g��o��s9L� ������#�����딑�	��dcf1)���s�,E mY�)D3�0̋^@5;+��'���_�.2�\�o��T�Ĳ��$��d��	l!�)�I�H���c��^uE�<#`��D�2	���E�8�d �B�$l/ےP�4ex"f�$�a@W�2s�q��%dӖ�z��O����
d2��L�nfհ5�k���=��:֭^����X�ݨ[�ۀ'F����f��S�cJ���+׵�X��sc������%�A�^�lz��$�c����lG��<���0�0��@�KY��5�1����5�ljkp�O��Ei�[[�2o�*���Kx�]�TR�1�

��Z�	�_�s�}
s��������������U(>J��0&�-+4���_Nt������(�Ѕ徆�NPh��r��"͸��J��Eԉت��R��Of[����r�Q"�akk�j4���=f��;�m�O11,X�����g#��j��[u�v1��Z2=���Av�������*;S�m��:�?�-�݌�x-�dRNք�G�����-����q<x~�Rv������g�y6i���O���?���%a�]������N����ۗ�e,�H�����
o�j,�"=��͚_s3�d1��a9�Z�����X&FJV�v�豣��Rh�ǎO_�+x�X�K��Y�N�Qp�1������IHm�*�k�C\�����Ξ	�x=;ި��dz�����$j��h^�{�o\�����)�>U�ۥ	�XH\���\�2�aQLƛ�5[(���M*��M��ܖ_@��Ğ阅�p����H���z8��6x4dfZ��%@�$�)eR�g��wCd5u�زYˀ �s��ضذV	��G'a@����ф�x�?�+ /z$?�>�<�Ͻ�s���K�2�oh��"���y�ER�ߋ�Z&�PN;���Σ;^��������<�oV�h��H�ZZ�TS�Eb �9��խլ0
���������q����c~ U,x �5�$��$Km�����6e�,��h�����5��yf1j�&_FBP��b&�eX�p�f�I3KK�	��n+5��|w
�&CU��YP����}�S6���p���0*�O�-�+�[2�hs���+.�N+�sa,M����?	\�f�QO������q�<�x��a�&��L8Ώ5�/!3�l<�V$(�G�sD&sM�[�Z�km�R��V�ls��~ǖ�vC�}������{IŲ��ҾyL��q�6I ϩ$����nX���st�(B�qV�)!>�b?���d� �~�>�v�2 |�c�����m�i�Y��9B�Ɲ��nn�¯%���5���Z������k�;�<�J���L)K�4~V{�t���0!�av�VY6t"�D���(|3���0�������e3;˿�Su�<�/��n����;����o,)�	5�صP��W�?\t��p���DX���׌!&v�N�+��;M$�4�1;���+o�(����k��>�܇�/~��D/\�X���ߔ�_��pW���<z ��6���㸆�d74;4�bz���:�	�I%��"�4Cj\��Y���>�\~6���Nغ]�}�K[��:%4S�d�����Ev��2�׆�ԗ���l2�gjd���5���1(��9�5�(�E@hz����.������PQ�����8a|Y ˄+���j�G=�f��7�^��m�J���tYt��2,��Ap�yjL`�ɂ�j��hPd���]�f�Id�ʚ��)���5a4�k�}�)�G�1�>���q��5W5=>ð��T�kC��5�͖s�IQ_���v�,g	�vn�!����}��җ�½�V��/��goT�t�6k��ʸm�B�S�N�&a��d e�"��������3�]�_[�vs� �p��-��Z�����Ci��*l���VM�s�,��k��y���AL��y�d�,��� �kC��0~F�8��(w��q�
:���hKY�}�;���$cȹ �.�	a��4i>S3����2�d��|��1�k�0�'�"̲����-��CV��6�]�2Y��Jc,�FѹQ�s3�y�v���m,���0���f4��P�!��}����x����k�1�AK+<�&������w�o�U���-��20&^��kȝ�	~q�Y_�ι�L.����*a��^>�t*���Q��D����������_�g�]%1�p~���^YG���E��qk��0��11aI~�������$��ZЋbfA��F�:���y�9 �u��+*N�@&<����Jz��^��D	�Ɇ����;��n�/�,ʠj2�~YS��/:����lԲE]5
lö?��~\���3�bV�x�*េ����C�$N��M�d�٭�l�<�L�X�Ʀa�����k�W�����g�Y���|���7����{�H>+��3g��I�������ڣ��}9Q�3�F�N�օ���G�Qè�S���B���ZB�^&�ſ�]�`�=G�ɮ�ݾw����lx��{��6-�$"�I��f(��eюIi���#H�F�"�K����taqd6���̎�g�0t���sD���\v�v=s0�ca���v	p�&��"�]9���2q6�(>F�:4XT# ht�@+�p�Ȫ⹪�*}�ݽ`e��E��.�>������0g	����*Հ��R�5�(�Y�4�=Z�.j��K(d�{Y&-]Gq�v��+���6��4��ئ������<��p�L��Ic�>�h����������?�Gա{�E�v�������[(n� ��:�0���
\$S��W�@p��#�޿�S/��u� �����v���$t�^�<;+���0%�$(a��ѻ�lI�r���q�����%�!TC(T���E���Cџ�&#�#	/-�Rh�
�`�YNlǒ�$���;b�c^�z+ϫ���M�j����f&A=��!���۲�Z�������s �v���{ �f�H��<� ���@ǍL&�0�~%��v�k3R������� �Y���J
���j�WI�2�дO�e2��s�X1x�7����f��(�݌���2��s2s�{_����&p�=�3�d����̝%Y�ٲ�,�
i�빴wͼ�@$�o��@�~��v���Zz�{��ٖ�3Q�y1��\/z��� F\r�@~���N}�,1������Hgw!�v�-2FE�:T\#,�{Б��?�k��d��lU�Ne�`�.��m(��Y�_~�m-�~Y8����]W���
.aA�;#'v�]e��� �.F�O�^J����N�|v����IfLv3��>�Y���%j5}��>S}䓟ů����ϩ��:��a��=L>���Q�c悐m8�rm����:�,�����$��Xe�\؝�5\ta��],x�([�݅�P�o���fY]%Ŕ?��#	�������k�r����Fg�������~ݘ�	JzX|b)��K)J;�ٙ3��︳]�ZL�/u�J"��#ì6��T��}WR��s�j��O{,p=�9ګ��x�7i���������I(NsIC|t��H��cA�e��N�z	�
@#���z��q�,c!#�oI�����˚�g�s�'
Q?ٖe�X ��iW|��Y}�n z��}d�E�2uh2�j������)~MD�/����G�goN��u��h���� ��hg,h�ܰ�e
k�v5`)��"�^ ��j ���M�v�tta�y;D�2�
�ȣ1���?�b����+�l�!)`H�n��>�.k�>���E� ��ZX�.A���u��eG�|�z���
�X�6��g��n���ֹ���[��m�����+Xt�;1>J��������Y�&QF�_��Q|���!)�]�^e�W�z��x{���Z��tƶ�)͢N(��Џ	���*�0�%�4��i�f�1WhU!xL�x�p�&�~
"ݸ�
�M���?m���)��_�v<T����Y�+`����)�oz@X!�\��~��9V���l���LL� �,*,f��(sO�Y���e��
����}o�;�ySה����SS�� �N��uM�O�i'��3�`��U�z'� ��z���o���N�oR�3�
���W��PO6+�n��n3hw�I��"�.n�I��n�Њ@�\����T{���i�,��Ggı��q����ﭑ.�A;,Ú�|�Bu����#O=Z�/��P�o���]���տ�~��V���7R����Jh�@DA��c��.�I��0���4e'^Y�!���0��9��,��Qf1�b����:��s���}���ԜQ�\?�����G1���w~���.]������W�<���@��E<46;i�����o�)��Hѻ�t*S���%CW�J|>>'�D2>yF2\f�$e��u�SWP$�M@a����?"�)��8�ҟ�@�iw�o[y��d;
�=ݣ����P�g\j��#%���~��)�����~ϽO&���:\T�&>oǊܪ�2�G�����4�x�u��{�	��?F��ƪ����:\}��_���������_�ߪ���"~Ɣ!����B^ec@�Ȏ�e9*��ֹ�:$26��cB=�,@[�ע�A[35��8�w�Ъ�b���}�y��/[�脍(�e�)���S �U\�7��l2� ��x-�krr�q=�Bb���H\����|j[f'g��º�U�ؒ.�I��������31I!Y`�"	�1��l�ٓ�th�^{���Mˊ� 4�0��^=�`�-��Z#�>y� 5dk�
_T9�)S��ܶ�P��jF݊L��� 5l5Y���k��Z�9��j�h��<7�j1�u��`eO=/� Xy�E�c��\˭~� �[��L����<]c�[,PH�?<����m������ ���5���x��FZ�͸n�����*���~i���Ͽ��c@���0 �e����RDyb��0�.%�%�ă�]E%;��gg����֎�<��]@I��pWڼn�>��k�N���G���ɛ�P�]\5;8ź��3�ze��d�(���[��o;�}'W�N���	y�/�y���㿨~󋟩��_���}	�]�4��縮�ս�ӻS5�W����ݻ'�ڲ0s5�9���؂��L�N؆Kה�E��[��ݻeav A2-��e[�03˨�P��vhU��t��	��w�P�<K����*�Hi����|%5�.�T��iaR���,�yc���`�6h��E{�\��
4b���r�2C�R��d�	H]��'��̈́7J6P2M:>s�m;6~�z��M�s�ID{	ɴ2S���s�j%[�s��/i^;�mY
_9/��Y{ �����~,�y������X�&�v+ud
�cO�p�!�#�t�2��*5�d�a��a�y��,.]�Su �F�y�{8���şV?y�D�S�0\'�����+�՜Rm� 6k�ύ��(�ER���΁d|VQ�m����O�GF��O�4����h�W��( ���Q17P=[R�9�B\۠���]��h����rxr��"�6���>2�BJ��[Ԋ���q�oē�0�ď�Hrg2�\�K ���,. ����`�9N"�����y�af���=8G�Z��p� 3�$%��v�LN��U��ϞO�1��|r��&Q�l>�F��0?�3�跸/5��8ڞ�N��{��R���Kvt\�����f�X6���s���O�QT�;��r�̅e~m���X�	�������l<�gkt�w�ͷO\����3?��HF���<�\��lAm��z��;������d��A��/t	 H�^<64�rF���� ��Y�I`6��8��d�w˻����	�	h|�	g�*�P�`w�̲���W~�@�wR�ǅ��%�H-�](�Sg�\��w�p(����@n�:�C7>.xp�h&����)�|g�|w�?����^�J���>��S��_�)�j���~�:s�d��O�x�����/mctx=���;�N��)\8��(��m֕���A�ZN���<H��s��;�*�Z�42E���$Ĳ��ӗ*΄�]�
����9�e&`l2�Wa<�s��c	��&f��鿛tv���6�h��BY��ڑ� ]@e�ܥ��š��
K����wQ&��̳��K!F�_ّ�LɦI�� 3nO�45��f�����^��D�6�0~�VR;��ݾ���<�G
���~<~c^�	�`m`�s�.J���wAZ�e�nV"B_BC�d{EМG�.8��[����4��Y@+ |��_�Ct��"�������]��!%�� �#��0.�[�Mͷ��/�/Y@�c�覝���o�/�5R�b�q�S��9��PT+�J�׵r!���l�N����+[ŝ��!&�k]���1C`��;	kLB�(���c����l�a7�aDS�Wn"v�ωw�̭���F�BY� .�wk��z��9��1���)@h�0�F��K�����yi�i�.��h]ʕ�v��i����{�@��K^��,C�nR6h�ο��wY���,�3�2�̿y�֓���G1~��u苹y "sD'�U�lf�"�D�N<w���W�����0P'�]q��ǒN횩�<�H�ƈк�~S��O�9F�n덧�а�}±�l���&�`��ز�,��҂&,lENЈ��~lf�e��׷E׷��{5+�3�&x��n���+��Ǧ�]��
9y�������Y@���l���+���`�g��#;Jw:d�O���0$���b�, h'�)㧄0�ih���-����O����iԝ *L�H�	qg���<L�e�s���JҮ��0'O��4�b~Z��Yteڙ���Y�-!�"|ܲ0+��oc�4>_�ۿ�V����W���/T�<�T�ē��L���Sb�G	CY�t��UH]�I���:Y ܝ{��B� ��L����q\�|�bv�f�$ŗ�4E�˽���eA{�ĉT�w��S)�(��Q�����\�k^��v�3:�;5r��E�����ڰQ5����(@�!}���	�I\�gd�x2�"�΢�+l+�.�����Q���)^�l���Ze>�[P̟
\m����Jh�	��{�u�Y4e��W�w�O<�x���j�n�ݬZ����S��얟��V	�(tm�B�52�;a
��9y�,�]��b�V.�-U�(�j�ϸ�7���~:M��	0���M鋏}Ⓞ[׫o|�G՟���Ȋ��.����mC�ҹRM��Լf��b���e_,�<�.@���ET��:�${q��F�&�&�2{&�f֖E��y�l���`��J��;տՄM����@�]~�અ��˳?b�8�5����X�	�����a�2��P�b]�!H�x@^A��m�x�"�_��V[�i�k�玙�I ۦWSxk7E�yH ���\-��^[���� � �!����
x�p)�2'��;��h�m@b�ɶJ{�{ۥc�v Yٯ�}���l0Y��ږ�DJX���[�>���P��w@T�Q���>`
�H��l�.u��N��2CxN�ٿ�1�����K(MMVQ�o����̧;��z����8������yZ֯�~q~�9�ߞ�o���F;���k&�r����V�\���@���������D����1�XqҴ�L�ٕ'㣀��C�L��v��B3��5եˠiv����ʎ���|�����61�۟k~�sǑ!tњ4�#',u� aw�2�,���eL�tW�P��g�ً"���\����#�����ϻ�I����	4#��g�O�Sq\�	Z�W^y5� ��;��;ոl���{	��g7��Y�X@�;^3Ȗp��  t�
ÑZj��XWjI�9�}`S;ӜYdwq��U� 6	X�tq�A�Lv��Oօ,tu9�&�x�h ǹ,* ��H�'�h�U�W�Ҹ�ޤ��u@�}Ȑ�����!N�~OP�ژ�	-���D��lF�+��AX�.vㆭ���~�{��ޓ�����.��l����}K�-�#��?���`����֗�>�����#�!dJ����5ԝ�n��&-_!��a�{�C�e�K`9���6	0ǟ< �~~���9�����3��,f���i�淿[�s�<6�z�U�C֚rg���1�9�`+d�">7Dh��4��x	 I��
|�u��)!H%�t�cT��nʪ @�S������3�If-� ��[�K�q/@`	1���X��}ȔtE��9Lê-گ�X�Z:�F��M��%�2d���v��t����Lt�$����nmy I�K�>�K<+X%`f�@���{���P��6-��fd��l8�2�/f�]�vP���n���n� Pl��ɫ@p��oa∆V�/���Li��\�:���<=	�T6�dt��I��J��;�Z� ef�	�2�r���Y1��4C=LP|��Y�z�5?�d�=c���9�oS0�Z@���&�al��K��̱;W��7K�6�;��{�6o��~y�����c@P��q?u��O|�i� �b?��1D1�*�E���7ġ#��L�1,�;rctXlD�LX�H�E�v���uX��%t&ع=�n����Q�Xv�Iv���peb��k��2�+Nf��5c���.
R�HR��qפ��� �\�3��,"�sj{ݸ?��䪐4ޯɈQ��̄<�.TW�U&Υ�����%�Q=��C՞ߤ���d�|�J�7������?�1��r��_����;��n�p�͛ �W������KhXȢ������Y���v��'m8Â<K���Ñ�G3��-L�h�x����aZ/�ݨ��O?�Xu��u~?���s���_�������1g�bg<�F���+��#ۆO�9����\��v���!Y�"a1X$esd�4tܞ���"���AmjM�^D�.&2&�8xn�dL;��e���(50��A���Y�{Y(bՉ����a@ڹ�I�8�{bJjyW5K�n�m�:|�q�p:�@.p�QL��G�S�Ǹ�U���=�����ڻw�Oㄅf#h��/8.�QR���u
7s�0�9x�`��T��w/�C�Տ~���O��~�*�G�����r(�e_�h\��1�y�
�-X1{�,*S74�a!_��Op}3:`[��҅;�ұ� [fLF���2֗�ڤ�[4�/�p�,���&�2�v,��bY����"ژ�9k���-��q�[�Y�cr���0OƓ�{�Yd�� 7g9?�\5,_�4��.ѧ�xD���SS2S0X\(�Y��[�&�ː8}K��cip�̰Ycl��ء$�$���[���;A})a\���9mF���9L��p�p��cq��ޠ����n�	��D�R������(c�u=�am̘$,�y�AB\_�N���(�p+��,���{��斲�`,���ۘ�&k�>D���#�_6-���V�6�(ګ�o'�dN���S���B�6� 2� ��<]Z�BR�e+
��r����lR�[��w�Ӈ���ڭX����p��Ăױ�����h�(XG���sLS�s�atR��0أ��U�"(��ĐeU2$�MثAZv
����3d��EjX���ڙy�q;��U5:��S��&M�d,J�F�	�]t��/0	-�'cSdG�h��n�X�2��RsGY��ӗD����	�.�hV�X<νw��w����3TZG��~��ȧ>W}��_�^��OS�ݴ��}��I���:K�py`hڞE�w#�\�U���^�V\������s�;��a��uR��6s��w�R�S]�Z��p!6�&���S��:�������l�z��D-�]q�rO�O���1�PRe �!��"���~��x�6v�j1�cec�������Ȃ=p2�4�"@kB���ނ"۹�J ��o�����
��ÂQ��hK8e�r�iS7���ǵ��/:�I:�,�$�#da	���%2._��~=�.�s:4u~f�E:��u��f(S��d�&�o�}
��ݰu���V��}��s\��Ç���կ�v��cG������~�굓�~��xV��h�RZ!�]41vX+�odq��� y�^���-�Br����e�L+�� �C�ts3�,L��c� �,M�^ ȥČ�f�������eֶR�+�GL=��棄5Ͱ(���(�����s�E���[�})@i�!l�Ȣc\��Q+�A�Ox�9�c%>�l~�H���(F\֢okP� �U�h�,D�KY�0fN{�����(:	XE�hj�sF�Ļ�?����%�FF�����j�2�$�B��9�>l�kd�ߙd�|b(�� ���qތ�^�"pE�ZCȄyU�����@N�� l�WI�
��>�_��E�Oɲ+��m-PN Oa��V�+,�ϵE��$���9L�C�5_�Ђ�Umt'N�!�:3w�5&��:p�<:5��FZwa���wbr�#�T(��<z ��tԺX����.-� ����m�tb��	me������� ���k� ��8��A�|vgȬy/���m�K|����[��,�.�n�zK� �������~�1�IJm�#%.0T�X�tv���%��b�!1Q v�jt0������3�6߬&�}>��S�W)x��#W��ַ�wϼ^�:�v�Q��s�Es�������N�ʜͤcƛ(�j��k����2K�	�	6!+w_N��;kQ�B��hC:f��1�� "ݨ�<��hZz�}�~x��{ki�B���K�g'��>Q͌ODG#@j���rH%M�g�!3�b��vJ®lϺ�Hut�"�7&zu��c%-��L���G* _�Z���n��>��c���^~%`F��kBhCk���~t^�c��(����ej���[��QسÄ�^�Sɦ��r-	j~c�($; s�J��w�l��"��ѽ��
�%0M�6O>�t��3O#�?�sY���kߨ���It8dR�l�U`rf��B�b��� +�[`_�1���؄~�{�iJ꺮�%���5�(�0�F���gaͦe5h� +��uq����YE�ƿ�`xԧ@ C�d�,�e�*SCa~�s\�p��y�,�!����O��i;��(棛.*�����U6���b<g\�� ��j�$t�V�v��9&s;W��\+���4�s1Í�v�x�I����
�:��z�"�%�~�Z��&�s.��d�����0��{b���$�����[e�ޔ|�+v���A���W�~�IR�9�̦���Gd���_]LZ>G��A�l
45�<#/���:�����=?7B�R6�8�}h�n���%�������B��*z�@;B�j�<�2@xݲF�F1h͌��T/"�t�����o�;1��Ȼ5u0q�R�&�F�>��7Am�����5�2s���ATc"�h��b���v�ݝ���eMϯz�;Y������m!-�,��2��1������X{��9Q,1 e}\����[�b�]����cQS�"R44�TW�}J��b�Sfݲc���<��X.�;9�������52���)�����O�󗞮~���Uo�u}�U �  a��x��������6I_�����sq��P���h�@J���TWHM7D�F5+�;z$���I����8�&��B`,�	�\�L�8��O<]��+���������]�x��&��ȉ�l'���r�7[�*�hv��,P�q��7j~���>ISh�I�L��d~�?Sv�{i�y��3�c�N��Xp��}o�n>A�.~?�qG��*e3`�,&���׷wמ�S�a�bp�w<�k�����b���5��XulG8��p�ޢOM":.u���r��rSh�d��=����?p"�����:���O��E%>�1�1ëPc�^@����Y���ê�#۪�~p��n����9
�Α5�Ņz���~�m64�ոbv�AG2��Eڸ�Ynv��dN�x���d�2=��0 �h���������t��4����\�--b�)��2��ր�?õ-��%�ϖaL>��R$nF� �e6�y���a� Z0��,�"�,���4X!��s�셂�A����<AD/�d�vzs Dg6o�BQK���uDٲ0,�k�������8f׺��gyf�������ʒ�A�.���ϷR�a{����5���W�&�MsD'��ǵZ�L�ТsN��N2�4��v1�v܀Al@��L����s�	��פ?h�(���@�������Td9^
E#�_��S�|�39 �m���A���dp�G�j�X��/j<���"��9�ߚ�9u�i�fSY�]�U+5�ɯ�F��x@p�Z�����������_��f����1��=R���'f� �駧'�j�dЛ��B�����B����6m[ �/38͠�U���Y9���f5��d�u`٠`�ԂBJ�)T�F�23u�I�<��-�u�dL&Y,VI;U4jE�{�'Kh�ݾ�2���Ԣ�@cO[�����-�n�^-0�@ﱏ��:�X7��vv��gX(��'�K��V?fA}��G|��O��P��j��V���;ի���z��k�c�>U�@H�"�LVl7����c��J.��i��w��]H���	81�] ԏQ�<��8@̝V�~��1�D�\��
���� �FY`G��e��v�'�~E�#J}L�%={�ɱ�e�70����� ْ�b�0$%�PCqN�S_â��E*0�I�RL�Ux|y݂�Yʑ(X��M�X����z�0̞�|��N>��'s����|Q�`��b�x���(g}.���Z�]��nh�L�	��)�|�]����$Yd�ػ��cTu�.N\uVHp� �����ꓟ�tu��Ql&���a��oWW ��u�F7z"�K�ο½� ؞zߘ�-���g�Q���`��"�*���ݍy�J.�|w)�nO���@HQm'���c{-	k�u*� ̪^K!�$���=S�G�*m ̶��~���,���.�">����0�lE�I��;8��Iv�������M�䡞�  ^�IDATw��Ӂq�0�� ,'`���B�����w�Cy�^�Έ�\�l���> �(���C�n4l��6�9��}���v�Ɔ�� �^kxq�n�6��=Z�w� �o�:s3F:��ކK�M���c,�1ϥ%A�]Z)�ח!�A�V7d>S[�C �8'?m�N�������.6A�~�c���VW�f�:����Pk5��������	�A���znnB[��D���O��w��;��/��@����ؙ7=�}0�[L����1tz��A�Z`�ڹ�.��e��B���#@�3��:}+��0���,�0��)vn�H�~�:Y�F?Q�bI���2�J�/�Oy���<8~����L�O.�Ty���q�.tm�߻�w�C\)-=��ՃX�<���A��f��X�7uQU�ɮu�Ƃ&guɌ��`G�xP����"���:���mF �;'�_�E!�)"����@�0��]�q�~��3���������{�D��_�j����|���V/<�J�ͯ�:�� �5|$��ko,��`Zz�L���L��.�T"4]f���Ǝm�:!E�{��K��5R�,賆�`k����s��\�/����TX�{,0��6��Y���l�H(�~݋@JЕ����} �Є�&;��%��P:.��������?��hu� K��k�F��x���w		��}ݱ� ��l�]���LOD��TY<2�؃gՁ����2�j�0T浨���q�����.nW���4��A}#��'?�Q��'�ôS?l����U��_��=}��6I*=��@�Z�6K��-�֡[��(C��S��H�CV�"��!������l[�����EE�0 �,0?h����)^uk]��j5�2�{�f���@ 2�TÂF���Zi�8<���qn3�6,a�;펌?���-���eih�)ƏU�W�xd�Y-|�����s��紱	�cі	Xo'��
G��V(�*=bg�80�cM�L3˜�XP=�.	��dGBO�Z�ER@�A;���g�[fs|���	�l��-M��6��?o��m ����e��ה��9�UѸ�$-+Vaw,Yb�p=s+�&�U��1���4܅��+�8�{���ӆ��)��2!���{�Y��X�<V�	�'�Bp�P�g���$�� ��-�&�ID�(��-�����|�ljv��wJ�1��*r�{��<'����e��.�LO�񺎸}�eO"q�o�,�r׻X�}k�;ѹС�W�yE�_��Ѡ`�1�u���1�=�T5�s"�	��)����S����g�,r;���'�@����MM �گN_�]�@%�E/�H[���½���IS��Ǘ�sv$��?���ډb�35E{1�*a3o;��3i iBd��!'.�5����6���b胬���jb��_~�{�o�\}��T_��_��oV�<��O��W?��I�^� '@ؿ��E����~u����?~/�gu��y��ꩧ��ɘ#�/�� ��H�4ܧ6d�����
���/�x$��n�{v�r��)��˗/eR�O��"���{����)�#4�`��
��+	��������]�eY<���u�Lil&�����Eac��2�F0r7e���{��O�\�(����%��q	_��t"U�k��}+ETY� O~��y��O�w��؟�s�Lf�����F,���!��/��V]�|�z������V���ߩ��_I��y���Ͼ^��׿Q]�N�U�-���=�,R�/G���_리��fa��M��w�v3��~���pQ�%�ݐx�9��<���t&��g�����ppܧ��,��q�`HŚT3<�6ŷ�Aڬ��b��	�Xʹh�G���o���p�V�<S�C�ſ	��=8'L��{�j}5������֒�X�T� ����R��ȣ�5V��B�I�`�ꦛ�@C�2:�����RLpD�g��-\�(�Hx����[���/ox8f�7��4s��\�d�	��=��R����jwgS�O����s)�t?JU���gRO��d��%��s��@2lC̗�3�W�-d��c����R�W��(�5}��Ŕ7���n3 �"�[�9?�����F�̱;����&^��9���u2MYn�v�?͛�W�;�X�$�cK���\q�s\� �"��Ts��T��w_H� ��e�M2�k�;C�n��Ih	}�vQ�yH��@���Z�����A!F�i�_6;�ͯ
�5�o���]�Ya�O��;.�ר%t��5fi�0.{1�����á�)$)�,��i+-��H��g8�^��e�Mz���臊u�K�utBH��S���;j:�(��#ſ�=L fX{;��ⳗnV�}���oTO�5�������������Lv�{o�To�u����0˩���h>�#�{���r����i隬YR����eBN��"a늙2���a('rY��f�$}����d2�dTf`aR)��ｻ�'"�П�a֕�]C[�4��R�)@2l�"��"`HrvjomJx�О�����)��;{�0�_� ^<�$7�p�ڹ����CCs
�����R4V����� z�F@,�T�b�6��(�R�:�L@2H]��3\v-˙�����w��~뫿U=����1t^� �Sg�W����E�!�L�Q'~���>�P��A6b�5=Em�dCӲ�h� `o�'{�'�	A�v��p��cƝ	�'cj�~g�:m�(U{�A�����ƌ�x.ia�TX=�,���|���&�<⳰�����tD	t��$�BXR���m�q5EL���>Ą��)?$���|���(�X0����r_�åE��&8��]��R��#H�N2��:_&P�����j��Z`�d���k���R͜g~ETTM)����Cp����i!ǵ��]��cj]�Ϣxh�Zg�\�F����Q �C|����&�/��Q\m_Z�w�d�j;p� �C�t�!ع�6l��q����<[~ʆ���ş��v��_���}r�2��C��Σ�F��$���56T��Ty��4Ru�N�J�"�}��-pG� +��y54�zY��j?;#'d&�%�I(�����q�:~h!Si��K��&'��,�{�,��_;�N��_�[w�f��$5�.���;�/Wc��&|B��	d���$����o����Y	?09:Q����:�/6 �����u�s�P�e6(���UC��,�ˤD��}Hk�H1If�\_�%��P��x���?�T�j���kU�ًsh}~V��'�V�<qo��瞨>�܇��|������p#��F���u>�#G��X�._� �h��pf7��⡃��g�{����)�m��$�b)w���y�*\-pã ���/\�����E46��h�o�}�M.��C �ǐ���D�-Ea����v�����r��9hs³qSu��k�;ci�T�w7�=�P.�����x	��0��� �N�Uv�Meu�\��VA��؆�/� L�~Nf�� �#hS��8Q���O~��򗿔�(�$y�����3t�D����p�wWo�� ڑUBq.��G���e�k����F��b=�/���뒭��1;�{��q�����i��9��mP�ҥ�2����-ҷH�L�+�,��xvS�֕�R�!��0z��V���dE�k0Z�|���)�8�,�+�8���W@[�YP�+�a���&��`�M#��f�s�P��n,��v����* ���c,�fL1�X��$��Z6�]����շ��*��x��Ya6��z��9
��p���^�(a��ad�<��<�B;�E9�N�/8�c�FWF��Z7[I����,S�:u{6�:��@�ײ�jo�?eHU֮��F;�e.�FK��1���R[^�/s��m�]u0�A�.�2N^�b|}��͖�ʼ�����~f������6�QZT���}3�@�7��n�.ڌ�eގ����k@��ιj�zEH�MގW��Z�VP�m �+'��x�- ڐ��X� M,�R�|69k����ؘ,��V���O9���D"�`ǥ<q��)�z��AR�y��h�i�� ��lυ��S���Ia���6�{:L;��P�ˌ��R@�ď�sw��Hٶ��1���z�9���FI�9�"HD�$�Sk����R����}�d����U�\�;�U� �r���hں{k�g])'f3��ENl,h���r��'�]��#�	��N����N��{0�ŝ��l�����p4Hs�����U?Ǚ�^`�Oz�;d+M�O-�x� 鄻�h�&�V�,&8�n��� ���?~���kg�]0/��>Kj���O�1��r5�����S��o�N}���7^<�"�Y=�S�͋�v���{4˄�����	����H%�V�#K���6��� ��S=t�=���j�;,������Y4��'kLa��WW	a�x��E����8��xv���\h] �Z�Ӯe>\�]�:9���œ����y��ǝ�edl�SA���uD�t�M�k�.&�ذx�za}ܡ�����z���h�Ro
-ٻo�k�c��~�RL#')�b�!�>x�@u�
���:|�>�_] ��_����z���aH��>ڜ��E�Zz��U����և��'�]c�wɳ�;%z-]R<��Ш{��Q���R��a/����&�"
\�6ӣ�ؠtl��ٞ�6�<�����-�����Vٖk�Ds�6�A'�"!ԭt������M��ꖶ	��X=:���XP����ui��[��slv��5Bfz�M�z�6j� k��m������.~}X|��=�0�b��9���O�mF1�O���h)�u�25� ,�Tl�AJq�"��&�g<{����]�"��.�
��pZ짜�@��4�D�ѳqnk�u V2�Y@�����a��]楈W|���ޜ�j�HF��vpCՆ�����M�b��|���Nlr~���j[�*���;m�N2]u��v���E�]���H�����Y�S�m�Y��ݬ��,e�q��QU?G_	q݆�2�����CXFe�gO-���X�Cv^{��vIAa2M�w�j��B�a*�|�ZMΎS�V{a�:��V��ލN�s*�3o�Ѯ����6�>��#@��t�q(��2/�h�H��zG`�אm�	e�t߳WoV���W��H�ӗV�8�G��`�&ם����w�#���|�*�O�Y���M���9l%5T:�O�n�z �Y�\�e��"=�DȌ3H��0��T�]��ꄭ�3�N��5�E�u�P�r�g�X֤�����Y6�З���v)�i��U�^L�2F��X��i)�O���MŸ3���̗!�E��+�19$�`� �5k���#�T 7+F��5t7)��Ω�Շ>�z��{�z�COUOS�����Na�w��+���]�nһ�y�m@�u�Z�d�}�3��|��,F��~����܅+��.�������Ă��)���W�r���H�.b�G����<���g)���:�A#����t5�46����;|�BfP	 &��y,l�!�6ܕzG"r���g�/�wel�,J�`�d(K�#����jӺݤ��޻�:}�̛�y�M������J/]��q�A��y��L �Z�cǎU���g�/|��>��i����oW���B�ß��L�IsǱ`"g/�4]�>�����\|�Ӱ7f$)l׵�qd��8̌�v�qg��i�ٹ�dҿ\��Kj�h�v��%Td5[r����dX����.�=]�o�����ϺpKB��������i3��2�o�0�v|�"�[|O1�̎J�z~L�޶��e؋�ؙ�ã�y�qcx�kL�=�S;Yf��c̛�o8�LO%ȴǦ�������~J���y�F
����j嘝ۄQe;u�Gf�a�d�:���r��y���_����,��0?t�杺A� ]����y�x��BD&�ˌ6�O�X�>+Kc�T��2�����w���.�������~o�W�F�V�#5��Hj9�
�jFۦuC8�z#uF���A��AZː���j|6-�������泆9M�K�M����{3o�B�+���$s��o��9�7��&Ҩ���e|�3w�aN;�9�u
Ў/��P6����sK�p)��> �9�48�osz�������{�X��ǉU����u��+׫äXw�92L�Bńfq�F��Kh<��B��y�p�D�*å~�4��:f�x-���F-dvD� �1�d��Ύivn�:yn��4V��XT{X�&X�o�ђ���p�v�Ơn�X�գ����%&�ev���Ԯ�.�.LN¹�H���ܭ':VĦsL�-�췘l-+���Nz����F�Nd��g���˱#��!W�_�Jz�����3�jP����z��W��w������T_�U������9���Wcd���@�+窯}m����}'ڝO~��h�&�7�|���/S��L��C1kt�꧌�'>�Y���yaH�;�L�m��G��Sg�c߷�`5��� �ԡ�.�	�,:J�u� VE�����vMC_ˀ,لd��KS�l��A�6�Zb2fu�b6h��;-�{`�吵c�g�B���G3�Ku7�oA�2����t�	��v��4p�J�|��Gy����1�<�w�j��_�^{�M��:A1�vH��9(}k]:2�j�Y�����{��,���(��
��y�AB�������B3t��邛\�e�E�P�_�:K= �g�!Cj^1����7�4\x=������9N��g���U����.���_�K�F��9��&z6�6j3���BL,{�Ӆ���ƀ�Rn�����.L�eM,��h�$6�g��������Rö&�� |�I!���6����T���U��, ��q,E¼eX�W櫄G���&"��>��5]���S�^B�%�Q�S��l=��V>RD�F�`��[d�Y�E@`�o�	���N��E�\��Z!�;z)~ǿ�Y�#X����.�ư/�I�e�����u-�ri�;���a���J�Ǐ8��p�l�r��D%�ʓ�1��P��tˌH�����u����<W氥�Y\�W�D.�ʿj9�r���1,s�}�(��5�Y8���~���29a��Nl����h�J��M�~��#�d�}���=��Yb���j����e�fo�;Z���O��-:���r~���V�=�N �*`�coBM;��{bl��`n2��	�Nv�[Wg0H� i�*ڗ=d�P��%��Ha	.���*�b�2�SQ<j�v1̤����&H#�0Z'���\|d�l+�&���r�u*�[�p�(��Νl)Y`4�i��(�A6�L02/E����Yå�X� �k�|u����7N������W���V�?�L�q|i��\���4a��/V�18�y�Rꠙ��������z4 ��f�i���V����T��A�B�e���ݏ�M� =\-�v�52dQ�,���U#}���"�N��T�%4I���2�c�Q=BQ 4�⧘�������.^�P�Xp��'�!�n2�{�D��K/����6�|�Tum�̎��̹s%�	�!8��M��0�Mm��=�;�Q�������:~���H\�&���_��G�|n�G����p1��E�g]+.B�'Nʺu�T��Ɯ&I�lw��}L� q�
��S�[�/܄$_��d��r#�,�u7�����S�71��C r�t[���E,�����1D)#f��Q�~�PT^:U;]�c�Y�$q �+�M�P �ppjAE ���qdg��nLۚg��� ��7�*�b%%~�"c���yE��Z.�be��8Dll��!t�B�)�G���ٞ\׊�3u���9Fv��[y*��u39_l.`T|v���o��{_\�U��4�>v����2L.3i}6Ɯ�M@�%B̢LBF����oH���{5N
$�y�Wm���鴋w˵E�`�Z.(mj(x��~����$i��:�}ab��~��P�A�2ziE�|g_-��_~���/����-9! %�PlR�4�C���əbsry|�zwb�z����g[�o)�<��j�4 �X����w�y�<}�E��j���S�o��Q�:&�kZ矽���cW_�反T���u"UQ��w�@�R�!�h�9�^�I2�eԕ��b��x|�CI�lQ�䄀��*z����������g���A؈]�q  ���m��u��R�1ta TcH�X��5D�U��>7�Ên�25����I�����Re��V���E�&�uV;rE�}}CL�L��渇���'�=rh�C�"����&��,�<�0e��=鎬+m?�o}��hëק 2K,����q���a4D��[=����=F��+׮$�b-žj���Rߣ�e��hΫ��E��J/�C0b��Z��1����>����U=�YS7r���T��bo6����O1��[�+X�͘�K���]��a�)M,��(�q�s ��a��z�o|�I=7S���v&J5�s޷�}+k 0�a�b�I��wf�M��2}_�����GqXV���SO�g��ṷ<�Pahh\j��A���
.�+��l�"����t6{i�uU�%��U{��@3sb[��`��X7nb��X���4��MS��2+2,��]�Dı%��5@T����q��O���XCL�ӌ5{��Q�.��ݼ���&� ��w�o�m�m��~4����Kp�ކ����e\LêZbC�H'���6�$! �f^2���nޟ�U\���b��� �+��"�nYT��h�e����Xg:)��O/nh���NƏ�}��k����C�!�(t;p��@0�OM�� �ǫ�Q��c�X�q�o���� ����4��v���߈�6����6�!]�!�s����o�y��
>F�*YK��2;�	s�hv�P�~�gٔ�+ڙ ;�P[�FA�:=7Xs\�a�6�><[7>kn�t�)cв7�[�c;��j<��h�:��n�
��)�Fd�-��>�U=��V��
��53k���Ӊ�WI�/����O3o�sv֊� ���,]S��"k pϭW�nNU�S�&f���檫�ʖ�F�&!G0i(M.A�-1�R����h�;�ȑ6�'[�<�b/���VT��wͺ�E�7�.|��X�2�(��s�R�g7�%�>O�*�G�
c�E�� ���_;6M��m�PaA��dP9��j8�g&����\���N9��؁�j�P'%(.R�a,��b����&7�fv����ع�5�ĚA#d��F����Z鎐�-S0Hp��8],x�,B+#�(F�T�P}�2J.�Cd���sfb���b��*v�P6]IwU���f� 3i��;5�� �6������
���p�e\���_z�I4MJ��ބ��ۋ�б��>q�q��Ɇ�-o�M$�4� N�2�����3:�7��6+ExiƖmw���������)w��޿���U'�?5�������0� hv�� �cG���$��_JS�.�2c�)�bj��:(:���&n�2)�Q'L!� �gs��_c�� �k\bq�z�}�K���؞y�Y����:Z�x�����s�/V?{��B�7R�P	�_u���0�hv�,8�o��'4�'Lg��# l���v�aB�5D�Ça�!��`Z�1۠F�	 ~��:�V��U�'��};�qV���Z�E��R,,Ӣ��ks� p!�=c`]�����>�5Um�I����Z0^W`�,� �Н�mhi�l<O7��E�yS h��Խz`� ���"�tt_�*a �(�p ���}up�e��*x��6x� TW�tzCZ��h����z-�x��-3(��t[��-BG6�!�΃0��0K%���͟Z>�,� �U�^gӶU�KF����^��7)
VԥP��^B�[�CC6�|��6��H��O� 3��{dl�N,��R��B\;8+m�?P�N�h�6�#C�U�L�U�S�6з�q-d	C�,T������`��M�8�:��� (C�����V�<@�4���y�:��=c0A-�=����,E�b��9W6��(��:B�lZoG��U�X�z�ơd��{�d���ԍ��5��)��%.~��nٔ"��{�Dݠ����D�]DLw_�{� HA&#9�[�k����N5�x��%$��S��_��!C��e'8[}���ձ],lDő�a��Vx����q�Ö�D[.���<����- *���U����)!����9hs'��z�}�۰����k��c1��l��ʂȤ�tk�Y�*��"]��*�E�b�fK��γ������$C��g�����\|�M��א�֠��K�����"d�N���q��e��e5|%8�$�V�̏
d_jh��q�93�I!��܇�����_���B��@�P�s�&�y��X�cI�^��&l����<KZ�$,�@E��4�	Js�Ft�V?�鏲��.\x/!��#��җ�����4h��뺄��:u��a�����Z>�6i���^�!��D���-V
��~������K8�2���|�hv8�8~�S�JJ��K��s<���k�Kž��ً��%Cp��s��z�qx�ӧ��o��"� lۛi&{8o�NE���Ρ��5�'+�<[��uh��t�0Ұ���YJ_��~YP�Ҭ�%l��:��֎��<�"��$�1T��(�t�*���8�E����Ӡ��]������:a3F���K��!� �W	�U@��.à`۟R�xqY�B5h]܃�y~ϴxC�9?��LL���e2�d�x]�eVj�ҡ�$k��ȏ�|�.pAެ�׎$�T����֍������O�)������n�zDe�9�d�Ux�"��`��k! k��S0�	H��)a˵ �;(��@ǵiU�N_L:�K�@ky���G���"�|Wݐ��:1����aF������^�'�9W;� ��i�I���r�q/��i�`�UK�H��^β!�Bo�eZR�X3�%��2;5��WJ�(�5���2�y_sh�ƙ.M�Voݘ��$;�"L�, 0G�A\���u5+-�W���8(1Ȼ��������w[��ܿ����o~~���W����-20"3DѼڅR9X�ځ��,w�I���{@������(��}Ǡĭm�p��:���1o)g'����ZV�P���j�ȉ߰��J���+�{�"z|�p��q�r��A&���V{��4vfh�f2QC��S�hj��6�Q���/�,�~3��]�H�@-���&�I�T]'Y3�t�]�:8]Z4��Tr�T�MI^�'gc�o&5'M�b��d'X*[��[������Ʋ� �I���f�
�$��R �w��_0�����sY�^&g�����;�S�,㵇4�]�a
�[ݵs��ɲ8�l�L��9@�U4W�ScD�g�"��E�\���&I]�~�ӆ/�� /���c���5��񹸠d�U��dj�)��E���g{���#��x�@�E�C�ё�=0x3��]��41C8��h7��$S��wZ
t�fo��+VH|���g	p�nþ���D.:NԚ�����Zm��˶0��ͺ_ܓ�	gҺ?���l�Z��\C7o�<�,�����2?f�v�K���y��\���R~FK��Z!쁆�y������0n�s�C<cf��;fҳ�/f����]��+��>�\6�&3�r	��Zt��Z��Y��~�X�Ph��l��,0�\<5Gj]�����o��%%2I�du�}����������F�y����ٳ�3 ��0�kV�[�l0�NN_#��uf�͊�����>-��Ā���_�z<��K-�`D1�z��P_D�u���H����1����O��-��O�W0J�#��2�&K8��2�q�����{ﰏ�:
c�K��5��g�@X%�K_ڷk�z����{V�����#�Ž�Vm�6HI��n�"��E��[2��}+ߵ/)�B'��M����Ɨ��Xu\w���4�C��#bnƻ7��ȡ����[}���o}�����>~����=���v����7΢�n���Z�BMi�q�0VӚbF;��,Tn�fG5e�vwch6O#Hު��Lz`��S��TU5Ee�YO*�:�/2@;�卉��s)r�:�V�pv��@���v��e�f19�����s2�A���m���#�I�W�!����Ev��,�
|��vp+V���7�e�Иl$��EV�M�V'i��g��m�c�̶"K�e���>� %�>�oJ1��BO$ژ�P�yN5ϖLs�Z�33v�ޙ�;��*���,�1�.���=x�P�]��9��@����<b��b��hI�����HZ�w�׃'�O��%R�u&V�ꢛ��S������"�_k��˷�Fe���(��%Hp���I9ئ=��!\�e�t��w�}��t?6�� ڠ����K����N��LaghKϘY&BG���J������q�@O5�5�O!��M�ZBWfPhA�����	˨��^Q.�s�c,�(�s���P��Z�R���oPK	;��-Ō�ċfL�җ��iX4_�`���1��A�H���̧*�`Zax�Y�Q�[��9Y�H���|-8������"��ܸ���|IP(8T��}٧p&ؗCo�d�U��c0�� �HR��Z�^�۹Ƥ�"�-`�c	>dUh�U�Ҽ�g�#ʘm�5-�2	-xfL
�\�����x���a1�=L�<M������1.M�t(b�x�d����`DO�1��R�Ca4�9}�lO2w:L�ˀ��,��m5�|�~�u�n'�v�Bd�hs�a�k��Ǐq������lA��/�eJ���۩��*�l  NH���K�f͍q݈�	�-R#���l"+:�g^)	Ĺ���e�(�rIl����2]��_��Í��ԛ ��U|�61�4�k�@$����fԦZ��I�S,ԕش��>��#�a�$�+�	�^k8$5�ݎ�]wpť�N({Jk�8p��`r6)��?A-��)P�!��>th����Ev�,X��H����S�9����d�H�����tq���8ǻNf�9D���q�u�$l��Q2�N]���-qGZD�E�'y�!�D�4�Xa��ٵ��4�j*�{����`P�_��V?�,g�g�lC�ؐ��w���a�ʉ�Y�����{��ή��ma��W��m/''�"�N�%�J�|��hЙY�%�):���&��ѡ��vap�����~����|��U�s7a|��+J��C04�I���cU��V�29�W�¤�N�߬>��sY��Rqg�d-�1j���?e�J��ڗ�NXm�̛��bO�����5i؛&S�tzŶ�o�}�M���h�韩��o�O�s���������<�$�"����?�8p���p��wCm�*��[��e�΢�b$�ao�;�B�}%5���<8���\�ϵ�D͊)��$j�����j������G6��p��7kɄf���8�����r�O�O�v�j�E�s��쭅��;b� ��i�U��8�x��S��M��[PP�4\Y��lCR	�7!/�ӕc_��>��ݷ,�Q���MY��A��x����wŸ�v(�%c����t�.����о�q��6s����c=��"���*�N�+�]f'� g2]_�\�P�,%�_�e�l!�*��9|n�xl$ܬ����}Y2������Gd��-��y<]� ]�x+����Vu���j�ycX,\AOxK����T#����2�&��L����-Si[�&J&���� r��1�n��X�}m�:Mv�M��Mp_f%n�A�d;������9-+Cn:bA� ��ˇ�?�I���}o�;
e�ni���h^Wgw���?c�-��薁ۘh�����3C��ggxci
�����ũj����x?;�,�XhG`#���H�2&�?��C3���71���U�q�^X���Ţq3ԍ�؞����>�2ƫ�3f8]��P��}n�x��<�m;���rvɒT��$�u0f�+a��-���qO5��s�i�6�q�.Vͫ�-a.~&�.o��5�^�U&�Z	�I��V/$��s��8�g��0
�m%�"Ϩ�~�&L��L���7�B��2|3�nAq��� ��������e4Lz������9���"�ùϋ�jAO�9��!+� "@Ur��Lv�=�W�d�q+fX5Z���r�
��@�_���u
s:WW/&|!�gCYU�K0ҍ^GhfL.tI��lv�W	�]F�}Q���C}��WjAiTp���2
�K-�[��y�bV5
d]�v����0�@R�A�A���T�J�O�����C֥t��������!���\�����$�0�������*��� �@]�2���,��l�qC�d��9ZN�;Q�$#V��Y����6	x��_��PJd��o�r�m�;v;v2Xnv�^��3�ɽ�M���eܹ�q>��I��Y�oB�	tЄp��\R:��]h�U3KɊҷ�6h��q��IL�a	嘱%�$�$Pv�X� ��[�۲��m����C�Y��$�z��t2}������l�)��⫂%��쐀�6����f�81���}�j�F��d6�X�Xޮ�΢�!���0.�8��7ܞ�	�Y
�V��fA��"�k�a�+l(.¦N2'O�O�nj�:���@nK7n���o�{@ka�����S��m `yW��������A)��Mz�d�QF��R���$_�A�d]O�55�%��v��g�����e&V�(֫��a�̎�	�x}X8OG]4d�8	)�Qy���֍֡%�Ƹ?�:��.T7I�F��?�"����j��b�e��{E�E{��Y6�x�e�	�]/yMu���+�bg0#�=P�1^��+o�/9Y��*�I��\g��W�~����N�k�V��\��_.9�m�i��s�w��S6���J��eBf3��k8�Z
'������>,��B��H`�vȴ�^Dî7��6�JrI^��X�e�Ǆ �2f�Yp�)z)�[�EM����{w�ӂ�����fjی.5>��*�
)��9�ؓ?�)2����u�^`�����<6�X=`Ĵy.�!Wd���aE�uew�]o�L�|J���?�>�U|]�@���<�<����`���+��{���4 �������^O<��k�rYt��ӆ���]i�u�l��f��9w9@���<G�*K�>w�ޚ�����B�ƶe�U�B҆-!]ُR���ۥ��-EF��R����X��q�����(a����*&��Rl%+�ߺ� ��G������3̌���ޛos�\�,Y�,�v>�� ��ɺn�j~����p?U"찥��J�5��O	�kn)3�w�`����	�����3o69��|��d�1�����W��r̄\��Ę�D�v��zI��n��2/�~��e56+SCt|C���-5"#�FH����U�uٞe\-&�f�^� ��c�djɠ:ɰ\�����[�����Pm�5���n��v������t��{g���{���[�56iN��f|�#��pRu�^&C��G�����M
�7S8V+u�2)���5��!����.��Lu�r��Z(����V[.���g���j�m-��Y��XL0�n'a���^PO��Kyx²�-�zrf:���߳��X���w3a�
�9������(�ʌ[�r�MX�K��^gͅ�o>X��]��W�X��<=eYH���s�&ϝ	�ݘ�N�kh���K�/��l��eCa�H9�K��Rׇ�����$���1᭡.�f
�s�WJ�ZANaײ��.�;|�,�O�5�w�l����L���!M,����1{^�E�Yf�qj�ݜ$��[��.w����q�6���u�E��5ey�`ӥkv�\����Wz�d� ����+LH�j~w���.�-��򻝯�:@�y���ی��,w����]8���J}�vT��s��p���>A����5��_� ��V�h�<˂�d�J(7O������������O�B����W�����i)�)�ekd�I���9%�]�es��}�(�׼�z�H� ��!�KQ�\3w��[Eܘ�y�ʷݝ�����l�������>������X	w.F9�W��|�W}/bt�~�&�۰�%��9��Ma�[��6
�+��o����zaq�y�N3�)�����1ߠ�1���Tg���{}��E�|���mr/���d��nmz����������bb��L�7������ Z��AI�d t�unww�n�lt�-c]n��0.�v�Lp�e�+�����d_�	p7��	A�Y�CSP��Y��5��O%���Nb�a���%��I�AӪ/N4�I�M��١�o��h��Pٹx$��D.E0��j������['�r{ ��%K8��2�f����8�H��\�b)���,@�-���zn��������w���.-�E�L6^+��M*�\�r���ݺ~.�ٙ2Q�.H	�-Ϡm�q1S"1��֩L��NJ�[hs���{	�)�v�2�[-�u�t6L��@�c\�ez�~��O��,b>�l��4��t�5�K��t�2�F���5����wN�q�Ť3��N�-x���ݙ�̮36� =!>�(�[��p�n�=��4f���E�޼W�s���KI~�</����<�<�Z��{.aX���bК~R���8~�]t�wrfCV���f(�-c��RZ_p�x���,u_����`JZƈ}�a.���z-���A��s��GK6UP^[B����6�,_1�|��w��sAn�sSv�96�ՀQ�܆iXIB��y�G���1�m��!��c��D�i�T����ހ�$G���V/��<����� m�\J�ع��Co2�@j}���t6)}4φ�c�|
�	��;�g��uz��&��߻q1S�Щ��	�sd�	���--���&��g���~��h>	��h,yvT��u�#�دGWݯʳ)�l�#��q�޶�� �[��W�;��2}��������Q���}�RE7z۶;֠<��58`�DR�R������&i��/w^�t���c�3���p�=_&�̷|��y[��ٙ�E��G��p�%�Q��͇#Ek�A3o�����Ҭ�����K
4k���%�Q&��A�B�$Y��I2Ω�MY$���5��	�d�(�Y&�h�h��H�`��wJ�{,!�2�����
�_BF���w�����"�rt3\�;(�5�Yg��
���9��M�/&h��A�B����Y����,v�߉Rdˮ/!2���a�g{�v�T:����g���/aP^�Cai��O�W��,zfɔt��o�H�f��T͎��4�,�uH�fnl��R���5C�0S��r�Mվ�ʃ*��+h��2u�I(�X�55;�5E����f�g�G&�3��s*3���[C3~e����O��x+,惦Sx��������Y��Ci��$O�6n~�e�>5x�Po���{��7߽�V_ش�9�u�q�^�s`Ț�)����@%�����N��ӌ��������; �pm�ڥjϖ��^!�jkUժM���Hmb�V�R{��R�"�Ŧf��H��J��y����s>�>��u��:HUjI��*���o�[�ZGs�`�x��j�3�mɶ��K����1S�-2�ۻ[��ڶXl�����	C�Ə��q�KYҾ�_��D0,�%����\��q�p��S����xo�{9~����Z�����SS��@��ъ\�u�[\���r�=��u7�ւ>qc�}�QKD����r��_$ґ��K���m_W�Z	�����Y��?�	�vc,�l��7�����K�U<}aXA�Fh�yd�K	t�=A��嶸���6z?O'��i���F҉C+��Q�(�+�g���S�ʶ�qt0�͠��F%�W��bf��oI��G�/�t6�&&�_�
�.�>��9�K�c���}�>��{S�T�:���JV�~�8q���~��>앰&�D����h��7��%�4b���"ij��,�O���E�֤g�Zb7-��ć�me�砿�{IyC������Mb�,S)E������!n���>_�˯
�d�أ(;D
Ir����'��ɸ2b�;��-	x��d��F����U�>.�'>����Z�A���ËnVi��q���bX��n�6��6v3nlLB~��6��>�Ư��l��	|0���m&���,�s�+�O�2����dc���
ڌ�u�c(�9�xT=�>x)�%��EWfX��z���dTr�#���YSj0vJ���/�,� �o��H�۶A~�/+~���\�V蟾b����A�y5J�w�Nq-��,^�m���r��d2Z����ʨ�h���7	�|�$��&'���O��m~r;K�����U�A8_���ny�G��Jq!�,�qz~���<��{Q��z�ԑm�!~b�qD��e�;�$�L��ʾ0-�h�C�S٣1(f�x��"�j�8�9����W�;����������h�{fg+����F�
�������=�/�X�#�l����J�Vjy�j�K�\9M��"�!�b۩�rC�HhQ,����)�����\�����즨n��	/��EO���&dU����/��(��+S����q���m$ Øs�-�0W����B\��-�|������"|�s�����4����j��ޤi�S���Ϯ���.~=�p�"��1��y���+>�Ov������:�o�h;�^(�mi�coO\�mՒ_�҄B����+��.^MLu�\�Z=�Q����o��4��6��ef'��:yR#qX�>?[4uL�4�&~�{�w�܁i�^@�y�`i_�Ad\'Zt�ZG����v��e��g��#��Nw$oV�����ܔ��R�K_�kQE6p������F�����ՎzOˮ�F�Bd��w����e�zbLE)��nP�ݽh蚔��<��d���C�kz�1P� ��F���7x�R[��peՇ5_��Ig�y�q9y�N��d����������J��~bF��Mwf�%o�U���t"�+,`�r���:N��#u�&Ť�I��ҷ�i���Y�c��=��]�a���_2ٻ��Q���fa\�7�`�i�j�����t�A��CS�5T�߄��/G�]e��?2���I�ǽ+j��?�ظj��/����6�T��ڧo�(�r�?\���]�Ozn���7�MhKH�J�d�w��M	y���Kۊ|X.u��_e"M�s\����r�A����QR�V�K�vk>��V�ш������d3�V`x������=u�Ma���S<��u�����'r=dH�0�R��tD6Y�.{���s�'�a�TV&3�`UJ�$�Q%�)������`�,ˤ<��&��ңh�:���ؠ{{.Nta��	�F�0}�����D���h�sp��8t&�C�&W{�2�ad��/S�qinW嗀�����FAtw6YF�@��֐�S��@J��R�V9�L?7��W��+]�
,杨��f)]�3�
��K���R��;�OB§��݂uծ;����C	x����jI�æz*�{j��Ù�Z�X9�F�˧�gO��4�|ZױHd�J�K�h�B������i^��Xċ�@�.�E�z����������.��7,�hv��<�����@ƞ���W򶧡Ӟ��`��}*�y�1��gt��փ1�g���V@�����P���yV�/�]�P<��1���RN��S����'ߨ^��|)�貤=8<"�)�($U�����$�Ӌ�n�����Ho��}b͈��1_2�EHR�$� �2[z���o�� ��H�((��1M��j8����`�hxOn��2p�	�����>�!�\4�Sx�f�U�=D�W����+؍J���ȝ	N�ǆ�E�@����9툨=M��N�����`J)'���XlE�2���}���r�U�$�^~P.�b8����C/��Tw?<�o�`�.�/�����8��3)�u]��i2_�A �O�b�����7���K�%m�ۖ�6��.z�Ų���Yd�~���?��ap����ƶx��?R�}�&��?}������ex��Qg�5�C2Uo�6�
$�s�cj:M����=(�˲+F��h�K�3�:��B��Gd���_��@Bj�/E$��8#�p��C[ �4��4��]�-,Ƹ�9$u�^�YV0Wޮ�b�Q~��K|&9f*N~��"<=��g�-�aih�G�I�se;�٭u�R?U���j�����u����_v�CN�/:�FPr����i"I�:d⺥�r�89��L���;�Lr��o��N�/�/���r��.pd-1�.����c�j�D�o�ԗ�tW,6X���;B|νI&�G~�%��Q���{z臁1�Н  @;{XIxӠw��-���J�����C��/�*EH��P&ߺ���
5as�z�ψ�s9j�^�gK�Qe�s\��3M�*�䅹���D���)"݅�J�������ϮP,��<�@�Zqw�U����l):xA}l�g���(�'
��W�n���Λ�����������0����'�L^�.�'(����*i�Q��U;�Z�o(ǖ��6�����vN#R�;RT���9�(����#��*��! ��m1�!������������r�k��VaB�%4���e#��z���c�؅Y4�؁b��k��|9ƹJ	�έ�������}O�{{��Wz=�^�5�^F���&>:��>+ !v���rl��-v���s�����&N������R
��)?�?V.­��4y����1Lm�D�3����Is��d�7+	��pd�vT�a���z�R3�@RԷK���ĮO�A������{��
fdr�DN~$� �x+^}Wg�ն�\��c����+��9q:v���	p�ݔ�N�ޙZu�K�Y�T:�%ɦS��QPx�Cx�IPf���_��2ik3E!��O\�Ӡ����[�%����rcY�+�Am�?j�04��$s�}|<K%���6��}���
�xï8�&�T�	r��4,^�{����Gv̌R�W\_�]�.[�"LҸ�0Ӫ�$����}I�(��9���4�wv���*\��mx�.:�z|�B�r	t���W�)\=��puL���3e���Ld%e���ڛ߶A3ִFӁ��f�,�!���<y�z�ί&䦛���Q<'��9s���;��ǆB]��@�!���ItV�W��A�
�̷�lHf@�����cC���g�ܽ���:F�Uw�[������g�#��+VP��'V�`�k��@]W+(�T�O��Ak ܘ<��$�q�WΙ8<\�n@�� E <�Z5�R'��'�LGB!��qK��ڜ*����%�S�%��X���]����f�̆��GUT�i�|ܩja� X�h<}h[�~�1a����'�?G��5�uL̾�)sJ�Ij��I��\��꺡m�ɦ����}5L���}U��^��G�V��	��C�*S�	�E�!��ǵ�Z�!ɕ<����#U�[%��AS<��U�����k�������SZX,���屮ࠝ/Y�x���/F}Z��	2Fߕ��B�4 ��>������fQ>KI�ԪR�n�PdM& �k5��v���ԋ�Ԫ��N抟sy2�V�/Gp���7��^�DI�i>�#-���T~s��v��W���r/,�V2"�:���6�Ba��6�b� ��aD�ҙ³C��UB���&�G d�nCN��w�oЅ�ǜ����?,�ջq�_�'�?������8O��}�01�t��*+�c�� o>���I�ЇW���u*�AhĖ�Ͱ�U~\��pp~�����Y1]�W��p�?����_��Ai������k.����+P�K�vekѫ�-إ�B�\����p�ƕ`��O�]L9�qW����h�gȽ.�@@�ߪe	S�S�n�����u#B~g)M5���]��R̮�RM�M�ڄ�&��-�zr����N�o���6�d�h�潻?pr@�3��d����MSw�\Q:�>��w�Ʀ~�0��]�^~���Jn��.=���Y�j%fۋb�v�,bK.h��W���~-��Hb���l��M�t�A��$� +��l�^�c��8���aυ|B��rGs�-�T��^�NI�r�m�B�䞑����%U��eh��bz���%�o���rV"��Й��.2t~�x�/,�N���~��3b-8��`�!o �/�kzj�47v���2�F̂/?���-��`w��p��Fn�/��n+s�o_2�)�!��B��!��d��'DD9�A&��+; ���hZ�d��X����d��iU��g���f��� � 3|hW�\�w���|�h�S�R̋�L�x��+��2q���+Xn�`��WX�D��~[�ݰ�D���L^
a
��w/�,,��|<�8��.�}�ֺ?T�0*xd�)��-���Z�2PB� ��WF�Ml�Y��y��0�4wr���B�b�~9�6N�����~�ٴ�����+�3�U;.�d֍HwN!x0��v�Q�].�]���8��8�~�x��{�N�ѿ{3b����S��wR"��������?���u���SED{9���?�L�H�Z�!�� PK   U�>T|p - �9 /   images/cdb0e0ab-4d76-4fa2-8457-7cb33d05bd01.png�eW\����и4� ���K��ݝ�!�����.�qw�Ƶq���s��g�g�/�몪9���]��)/'����)EA��&�r�
N^꫺����/s��<�@�^I;�$]����/m�Y�c�(�?����F��U��+�WV���֣_�H0�n��cmt����%�80��f�^�:�M�D��O��w���S�� �>엡�����_������ \���S޳� ���i��j��8Y��i�#Ǻ�D��h �U[=��um#'G�tA�U"�EB?��"_���?Z-:�+���}���`�%ִ,E�[6�ZU��3����ykF"��B�>��"�V���y�p	��R�2���B�ҁnR%�q����=�Y��Z�ͥ�2uF;==��J�T����2'�q��4';n�t�u�i�aӶ�D�D��6�H!�X�B0+��Le��y��3tr�P�ra�-
�OП�[����_���c���w�.4H���Ť���Bޅ���|Y��}n�ѡ��6���J�4\YY�{g���K�5-w"�ˊѻ����mVTR�NH���ܓ�v��zo�c��4���K���`�L�L�R���O��Xf��
�����x��u�4��~�ZM�B�sM��4
,{R�H�%;p��cT�U��:��.�+�RE��R��-s�v)+4����b28_k+<GO9y���ы��d�7���yJ���V�@q{�Z9���۸�r�~)ؕ��#��
Ǥ��R��c�3pLa��e�v�Q�����c�{��cZrK(*X�׃"�7�۹����Nw�\U�k��?��Wۑ1�(�0\��1�Moto#!�H�#�N�Ԥ�0�c�?��5��!�2�C�Ѡ^\���.��U�'l��hZ��d��hWبYVɧR \����H��\��;>�Dc���H-�z�l�L��d�g����!�^!�hۍ�_̗��R`Zf�Ef��rA�j���m�7��D��q��	jlm�j�籕���q,q�T')����ˎLAL���\�&K)xc���� 3%���&M�Nu	�זt�y���N�GY����m?6������AQ�9�+ٹ�p��+P��o^9����bH���o�aH/�S~]����k�����_h
�cZ��,�B
�n�_&�^gi>�+f��&(�Ft�HX*�U�o+�hn]��U�(��Ì�"�,t��:�4��_Y���6��W�Z��/�eID3<hf{�C<��[�y�G��Xkl�%e�ڗ���T�5���c��G*�l'ږ*��n��5z/���o�3N+k�s5Յ��sk��������RG\�
mR�[�VWm�WpdZg
�j�kuΦ�w���n^�)��Ǟ?�:5�Mt���7�>�5�e7�n��d^�?��2���^H ����~R��3���v��sdʜg�}�Y�	�;���~	����n,)��M��z��fͩV��W%bTuom�����ۚ��_3�0�5T6�]?���b���͓""�b:5��4��Ǘ�yZ���V���qq77�5��?�Y��+**n'��4=���0���+c�G�@������u>�]����e2}�ۺ[��R�i��m>ꄪUkēm�7Iuj7w�nY�V��/�6��<?�/�]F�����}�_��(���������}Z�6v�����sbօ_��k���`�NŐ�~���<��'�<w���{�Ռ%掚
��͗g��m[$�@c���Y�H^�M��<N(XGH߶7�����aY^�yYoV3��f�����1���M\]��s8�v�p��������o�k��ED���=0�ޯ�@
VY��%�^%�-�ui/��g�ܶ��ti�h�>���!C@�75���3�4�M����ͣ;���<p}����2��|��$���k�O2����:E���F8	�1���Jy4������ƛۚ��|�K��E8��w]���}R�ߤ���{F��r�'�y=�2醪bD��@խc,��7�Xr��(�`'� �JPk!�1U�Ȉ����}�4H� ��}+��CȪ禭���!QH��|e���U��ij���@=�q9~�W�T�boL�P��d���K\��R�~��߃fR?�vm  $NU�Z�c݌������J%����E��Y��0fl�l���ǵM�*n>x��p
3z.%B<~{+�QNÒA}E�g���=Fk;��$�Ų>sǛ�)Sw�wV�O�l�{?.�V�3įu���rcJ�Y�}XQ�Z@ߞ56�������9�.�����Z�˙n<��%5��������Y�S��x�7t������_�Y�x����|����f��0���:��6rU�1���wٮ�J����2+~��� �%��iЏ2x�b\L�T�_���vG	是
l�����y�p��΁.��.�G�aj�$L�&g	M�$$[]����%
Kɐ�%5[��Z
�+��Zٗgg�Vb���Y 8,�.���^�~~ϣ'��&���6�V��������;�W�la��^̓,���B~�+�ye�|R��Z�d	b$	���AG�͒[�p�Jס#.V���{U��hZ�.��D����!asmh&������%Bϋ6�[�gJn���)�˙A��X��Z��u��\T���ىI�?T́>ӓLD�����x�y���������ă�B<R��W��$�*���@O�k�Î-�1�礞%A��K_�>��e� IB��YP;N��;�x�������Y��1*������хPc$�|4t��awr�5���u��08�O4���|�ŝ:�8�A��Y?௔:n�j��z9��*����i9�K�m���ȴiU*��x�^�3�V7�O2HNZV���hf��_;�	�\�b��q ީi�B�8�������j�iD�磌�-�����v��3��*���Hhoj�Y4< ��Z��23^vQe$S��FD���v��`�{��CF������Y�@����]'�"�'�g̈́$��żA�Q@�7t��v�fi���OdL��В�������Uo��O�m��_ւ(��y&�����I�����״�E�lD�榃�7�j:|X�&X�ס�<+�j�#~�KdH�+Q}����&�����>�︔r�d�ɱ��u���&f�7"8����.����7
|/ -7+uf&�Q�T^*�8x�oY/b�	��;>X�]�c�}��I�*�f�o�~��?Ț'�X�S�#�Q�v�\J�`,r���o�,��~g!'W�N��JB�xG�#:_K��¨(�U��5<|<H��®�=����d���;\��ϙ-r��tM�N�C=e~�&�9o���ڿ)�)�Z~@)�M���ı3�/w�Okp�s�W),]N�v4u�f�I�)���*w6uA|�fڃ��z~_�[4ɥA��N ƍ���O2��I�Ͻ��r�Ο�H�Q��#���:���IN�����_��*#8'�l��F�I_���^�MR� �$��Q�v���߷��2����T�d3:���"���-\"�#� �V��Ƞ[���vM�a��mh4����ԿK���V��[�R�dD5��3���Q�~�旤�XA:��]�ge`�t��^J�O�!�մ7�߻ߜ����'=Q~S�8�[����yZ��]"$Rl,nrQN|W�D�){ۘZ�׳���WR�S%#9"�=����dh���)6]�rZs���O3B�[��X�
�8a%����T� ̚3�"zì�W([[J9���#>w���^4���k`@�P�r7P��NA��#�l%&$�፜� "Nk7:jB:S����ܱr-2���'+��!�����/79�!G�X�w��k��H4E\B�Jԑ�� ]�`-QQAB�n��������+-�l@��t������$y��?�£+0�ܝ��:�wS4�v�`Ȉw�����|FFFK�u����˩�u�4?~C7Z`A�Y������1�����+��>å��ɀ��W'�E	'+Y�L,�_��'�*�;JC�/�\����K��/wF�A{����/��t�wXp����R�ˁ�}�CLa��n&�>��&�/|b�MD�;<��2�P��-���K� �Va�ZU��R�lF�Z����ki�I��N�.��J�����hFOs��殧�;�����ɰ q����TgsD3.!��	��ѥ5N�N�$�n*����8Ry���N�o�Dx�Y�v�0娫Ӥ��_�(ș�۷o�yUS�ˡI�h�kLv��,�E����k�g��wO/kg;����t��|߇-��M͜�G4�j�\��{ff1�������.���Jt���NC?�>2�)*�CO�(�	��|����_l�F{G/��[��?��.��(CO�[;8�oZ7���ߏ4+#m�R<�n~$����H��J[����3�z�3�����H0Y�4Fk���������('���z��r�T������{�	�K�9�_E��6� v��Bzz�of�.�5��?�\�ME�i�:啈K�K�o_��i�Z
S{
�妗!t���0�fj��wT�%f^��}T�ƿ?8 �sC@��8��`����|v���(���vL�R�}}�<�j&����|��set7�d��{�1����}��gX��J7��Ķ8=vD�� @��~�r9: oӱ�
2�`4JT�|]�����lǙt�
22�#��B�w�&�YΉdK���;qa�K~��ț�nt��Y�eGz�J����ݚ�0����R~�"�b��6�f.;���{c*�v�Di��_Q�z�#C�NyE�Y�2s�-�:�ɑa3�GF� �ݷx�V%<�a>�f���7�0|�����*]���#EF��rCv�(7;�4-�z�e�J*+�aiw5n���D�+e#_X��N�{���hBr��}�˱�{�~��;lU�f�PJ�}J�J��U.��n��oj>�~�~?2n�y:X��}b�O�0`12�<�N~�3�Ȯ>�x�HIJY��XȆ�8�55���K%����Ϗ(Hdy����N���l/7� 	"��q�ř��p�Ҫ�Φ�U%��R!>��v�D��REd��}�b:k�!~ ]����R����y��E[��%�*�.�C�����/%���6B,
ab�Ff��V� �y׳#��@3���q�q2_|NV�[ �ecBQ���ǲ�!��Ω�7D�;]<��f'��[K�"NɆZB��g�:]8d�F��͗�:Ma7�UZ+y�jS|�^�bG3g�?^	;7��ݚa�4R~[mu�!:��pDw�0���]�a/=/N�9��� 
�w�����#B�����j���V�.C�L>�w��l��\� 	ᘪ�&�5�6.��`!M0�6tweU�`M���v�����VxP[Ã3,�u-?�"):�D=��e���!!�� ��� ����������$<���uN�+CT���7?i��-��%]R��V�E!�x��8#P���헱%��������~�G�)	���2��"�(s$D��=I�AK��o�@���[�{$
���#"����r���7��ޖv�dy���HYz�v�M[tW=Oq�������K�� u��	�|��,����`��Xp�V�JX�3Ȍ��ϴ���#,��j �i�[tH	w������To"����9B�Z�R�	�K�R��J�,R$3E�^�V��9*���^�q��l^��!��H���,C����Ғ��y�PR�����xA�ټM#$�V�h�泯�������~���:v8�LLL����������m�7�E�Q����j_\���;��z�pZ� %��DԂ	�[�s��/%Y�ԁ������3Aԇ�Ѩ_T�O%�Y�'m���;H�_�`55��z�<"@�V�u�&�(�Rh�ʒ�����f�e�e�����-9�פǓ��&�c��2ĭ�B#��8*�I�����K��&���7��Is�m��3������+h���'L� ��xF�-�8�'���qZ���������=���v�uwe����^g���:�����/f��z���g����w�] ��ɱ��bK�$���^��f���Z=�2�eH#�~�!��&i�7���T���]�<����/���5�#�@fU�0O�u�`�S;�����,�^��`f�G����7���B��/�\�w��U['%?�h���w���^X�P��>,�U95�����ͧ�;��6���A/� ᖣ��4�o%�hD忘��#W5�H���'�$�c2��,����O<�}��Ѥ���
.|G�^⭋�!��7�����Uue�<*�����[C�Q/rc)�t�
TW'�����Ľ��R!Kތ:���c��z
���n~�%o*��:}b�Sj�CV��7��00C����O�ѥm.�Y��7Y�x����4�[[(?��[k	�@b��k����H{j^g�D�a�F�4��&8����������{e�:�F���ԁu��y�TI	f��C܃re~v��>�G�0�F�RƧj��/�st��i'���J�ޛ�u�~� ��ؤz��oA
���!o��c����9��Z�γ�
�Y�C����_�Qv��3YK�r�[e.N�'&bE� ��|��^������@����E9�	��SvY��-ֹ >m�Zߔ�L��A��k{/K��|K��PÂ�u���p�P���X�s�z�{!
zkH�^~��d3�ƭ�Dl���呈< Ă�7T��!�?�.�w����K4��H��Yh���Ş��+��ȭ#-m�1�'%�����0H��lY1t��[
���������!̦0F5co%�&>��r����)){V�WF�*�
�3�Fq�<k�����E���������%V���m��#šx�
H��j)���{�-[���1�^wL��+#|��D"��{CÉz�˵��.�$�LZUa�x^�Zjٝ:r�Tv	����d9��<�퇛b1�4{�U��� !Fmj0�6�Md_E�j_�唷@����{Hʃ�zy$)���.���tŃ.�Q|Q�����IDu�����G_��VG2-:F��*��+j�>I	N�ĠS���\��is��q���S�zSC�5��n:kb�R��&F�+��1-�b�6�P��Q�2l�EEY~x�6X�g�#��O��]� I^ 1Eb+����q9�E��n����~e��.5L��d+�&ۚ�רG6_���l�~���y�׆�n���e�:��+���p-�I.+�a�����4�y�Mڂ.��p�QL�[���d��v�Wdv��L�5v��n��ļ�e ���:"m��A�c�ͷ��Pj�p҃Iե���J*y����� I���%�4n�t�W�x��u���Bҡ��!f�4}���<bo,f��w��x"r^�G���#z����BCӦ%6#1���jj:	�8(,Rz>�&�ۑ�]�*x���� ���t��CXleW��k���r6�1Z�Q

������i-5����C`�T�rP�����T�%!['�`����_��O�Y��O܂��������`1����bL��22i�e-�XSa������?��鉶9-7"K�HW;c�3Țz��]:�/(�nU�9CMNg�� ;:�(�����D8il̜�E;���ǁ���)��dgU4[��g7A�Z��]/>?
����8��mP�Cq���}����z���#[����IQ���26�I����ܘ�)�1�����>���e��g"���Qy�+�7��?b���W��������T�tW+��H����:����H�i&�Wl����5�3h�����54uq���-��������x/�j�<K1�/��J]m�0k�Ac�%n���&��2�-R܁�'���uV�6�Q��h�c���?�$�7���4�az�'G�-�DH��~f�k��c�'7����+-X
����DL�M�s����� O�m1�#}�CkkI���� yJ�X'�N@JЊ���,�&(#���a[�{m��*����Idw����̲C�>��!$���*DS9��RE\�=h����=�w�a����f��~'�?w�����3<wFϒ%N�Zi]F��h�Xx�J������q�`�!��:bĨkB�T�iz��_M��:��i�wi�X��ݰ�?�VON�D�E<V~�G�}����;Mr����C5�kӕ ����mbZ���qM���݈w�S"����e�(&2�Ύ*�Y�
4���P��}-��l��19�������~_B���T-�|��!%�:K���J�<��(����ɓ�]������S]W����؛��
N��P�_�D��1�JV�u�^�Տ#?�#���F8�@�.F�ι�p�mꡯ��S��΋��*��7`:�]���p��R�כ����s=��#��[�L�3���A�|tS�
y������dWd�eJZ�ю�K���G���A�w�Q�ϥ��y�����w@*cg�f+N���(��ZY��&#��sqT4�mHgY(��%����b�WC U��{Y}�(y�J�G�#���D�>K���Bà��~������lO(f��������N� �	�u�A9��֋]I�0��"���}$�V�@��C�lb�y���2(�qlo&�	*_s�О鴎" G:�/C�����.n)�@y�pް��z�*�d�?�#{�I;е�ؤE����dʜ��7c~�<��jq��d����y[��CC���a�z/k�폅��v:���k�^�I�n����;���)�::}���޻yS݉jw3��Y����ʰp]ŖP�ǑG�����4��A�}�"q��_NM�&8�<l$B�`5�fmv�y])�����Q/�2Dڕ������9:��sZi�՛`V�O��Ɲ�1 ���H��;����q��T�f����1y{D�a��j��oѵ��}Y�$�9�ľ?x�,0�?��L�i���}�"+�t�&e�:q�U[�Ih�(�Y|T�LkW�[�R�ȭf5�������ͦ����2@]����4^e2����o��PL�t-!�fM�����k���$V)2�Xg�/%�_����[M ۩L��ÅQ�5���ޔ����@���ENNӚ�T�4(��m�΅�'�`z\�KRBa]�]���c��T��Y�U4uJiVư�����FHy�SR�Y��^�t��ϲj��K���-�g
����3����It��rS�b4�=:D�>�3R&�e?���6�g�C:U���XM��x���ʹ�F�6M^���h&6̤q�8c�A�D���:��,o(��+x�����Ӳ�(ZdU^`�=�����GQ�P��zI�,7O�]��ؼ ]/�J�<����|�������XK���~5냓 ���șG��� ��w�<�&�w/��ե�ٺ��qZ�QOJY�[���s��׎}�E&���-r����<��E}���\��0�F|k���s��߫�<���ΡO{�*{�?�9z�hk:�"p{P���^Ԗ�aGz=Zzn�&q'<�_�NƜ�5�ο�5�?#o��\�$'�LE��0V��8jb��pOQ�k����n��=��X��ܨV�G�r���Tڶ{�Ni�{������
��u=��y7��A����!�����$iM:\)%��f�)��}��������·Ⱥ.�Fl���L{�כ	d�#�!�_�0!)L��T�d���x?�Z8�8�,W��+Y���]�jғ\oU��������ZԮ��� �����-EI���)}�E\Rk�G�~�ܸ�7Co�9���S�&E��w ��
�}"�[4
fsOq�4t-չƕ�W�B��1���~$�K�9�r��;(��Z����?x��9�ϘOx�<�=������D��İ�_�g?�h����� ��?ԁ�Q�qT�`13�ʬ�&��iI�EBm���>�nr.7#@��NU%��Lo�,��x�eǺ�&��D�j	t�@�3]~�mDŕ3ҽ+tP֑�QK~&����Q�n&ĤA��݌]:�x3:[y=HlnER�^��w�����њI:v��b(����@C��K<�(��B��0���)���ѿ���&��n�H��/��΀GCP���ݺ�]�3e��dc�(���i�l�Y�E�{fw����=*���{�IB�?�jK��e�i��w����t��а��W0�0S�x�ٮ��0k���5mȌZW"�i�CTE��ai��_�˰UIL[T-���2�}��`�*�kQ��$v���_�)h�����5B�;�ev�\�� ��y�����X�?�[�ۡ�� ��V�a��ݲK���w�SiZdӜUO��;��?���0���mԂ����tWv�
��E|�CJ}:�����;T��/^b3*�;����w!����gկU��9��V\I�p�n�Q����]7��p�hgM�^��#(�.i�\v��|�����Ts�W��]�OIH����3�T�P� �Q��ܜ�E�@�kR�)��8��hޫ��������4.��':�1�0�Pm�Ag�>�A[9�I�76���1�t��~�u��A�Q��R՚�_5(t9^t�Xh�jNj+ծ���}��f9���5bHa�&;w���h�"��xB��&K�g3@Z��d�:zڻ��ށ
~���E��l焜�#�Z�sY[��U40!�Y8#����T��i0�.�� �|��	��'4C���~��~+�����/�dtxQ\��8%/T���8
�C�#c�o���X�yͫ4���'*�\+�T$��j�E�eᇲ�s�0��Jn��J��K�k~�cT��?��z�V��-�׶�?��f=�d���Ď�I��l�h��ǩ5"�5G�O���V�i��K��ah��)�Bdk��5�b��C�?�<��-�-���F��һ6��v�VqҚ��<�^w�=��@�F�o("G}p��}��6C���?�?�"����G; �N^�Ӎ0��ٟ~W��q�s	� ��>�	�J��fu��4`b�&R�?��w	���\��Ê{z��MY���'&�N�/~�9�A���S��Q��$h��gG�FFٹ3���Z��������m�~t4_o)�1n���ӔIen~
1f�q^�dU9�F&x�0r\�H�}��
Uy�s�;'��~~�RqŦ2�8��1\�Gc�n�[�̼(+OL��2sJKk��u�إ�����V/�H�q6���M��@�!�Le�+IP���o s'ů���)�19އ㛖4��f'�O�g��=��`'�X���7���Gr��01�4�ф���I#q�~4�/���Ӕh�fL��Q��&{تLA�U+.�'���b����-b��v���/_�!��ޝ@���2v��l���~Vm�:t=9=���G%�x,���g
����D2��vR_�h^���&(����@���� ��n�p�������߶^^�`��˺��-~2��/�3�zy1��Í�G�	��.���8��J��-�����^�Y��S+#e���ҟ�����_m>�:C�Չ��:C��D��j�{6j�w,�z�D�w7��EH6D_��}\R�U'���#���%����� к�O��	O�?1�fȅ�!Ԛᛪ	�#u-�3�k�WZ��	�p
�[]M�}W�Z����2����}�pk�}	�տ�z�Z4�2�{�vP�4������ҏ���D��)��j�}����gm3���O_�KϬJt5MtY��s����n� �Փb���?�;-�D�)]�ܔ���&�KF�$1�X[�L��%i^2~�<������:����U�J�Ir�9��"��#��a~������(�X��\��r�a�͓�Ҷv,����է�dͿA���9�J������3A��%�P�u����uƹ�]@)M��.�3>)����[��L��~#d���X�C�<��p��Oyh%��Mr�P�2%_�,մJ)r��}�T��JB�6>d!y�/��n���h�ƴ�m!�U��6D����#�r�|?��?!ψtg�S��2�m}}z5��:ȼ�Ps���M�m�O���i��	�4����Q��:�
-�c�@��Cm���Ba��G��	(����7HK����-
$����{;�ĩ��`K�w2�KR�68)�_�ga�%q���C������q0@��[��*���EjL��e���!��9�v�)��_��w!��R���|_$@s�dG��:�!\�/)0(��pwW�d_!z	Vł[9qY����f�%�+z������/ -�X.{�z����/c�Qpw@:]�;��#���a�6b�^6o��.���7̯ZNO3=C�|�Nc���8$[ssАHJ櫐�A�,�N�����ȶg��#7�pP�[�/��J�+_�b��E�FT3���rs;)1e��Gʜ��&զ%r��i`V�?�CO����)�J��N`V������V�~`+poW���q�����'	�(���{3��l��/�bTr���!(��z�J)۠)����G�ڤ�tR������i�՝��E�����T����+��B�q��7m��i;��$�ߋo-��.w-���3z�_�QII���F��|A���m<B���V�x�+�؝���jYw��I��?�?�/n���w�-����D��tӂ�!�[�����~�Qgu^��"��������ѝ\ىMG!�1�Й�X�M!�h"����SM&b��E�j�<�Іb���V��'�q�/��"RH����(`����5�L�g����
�{�y�2��Xi�-A=��72�r���F8'H]���iƉhϳ�[�{��r�e�����7;:c�����&(�K���f/�leu�|>]-7�ѷ�n�Jr��kz�1�����堛҃.��Q�
�b3���m�um¢��Y�R���Itl*��c!`�����H���2�1��VQ���%;��=���0��i0"��/r�&�� �m��,���/kov7��C����	1xOs3h19˳�ٙ�B&)3K�#6���Xz7��k�?9���+/��M�b�Qv�!��>��C�;�p��@���� ��be(}L�l\�~�>�&Pe��i�I7C:���P�jQ����(Mʰ~�#͌�^N8�%+7�	��<���ȟj����ò�Z���*���l>��9�8����w��t���X���S?�P�@�כk�"$�g�(֮��Ƞ7+��e�'��޷g���L������\�F��J�y_"�B8;���O�������:�/x��K�Ut{����`���S��P,���B�샟Zш'B�:�T���{
bտc %9�R����7�6Q�, eTd~uhM�.v�1�MbV�2�@��3_3����Z�H����ZiW�	U'������b���>����Ȑ�="Q�0�֪
2�8�9��\�Km�׮0���m�k�m���I���k�������wLR�^3��%���I�+��º�t��Q҇��z?_��?kL;b�/9�����㌿e�"iX��_�EZ�#*U��\^"���(pUO�[z/dS|Ќ:��g˙ΐ�G����$\��ף��K��2�J'�XS�Z��Wn��ޯ/���Oxċ��a~��WAĢ`Y5n�3&g��k�p�.*�o��\��_��S��/�)����w�yq��jd�0���΢��}�a��VҒ�����|�i�\�ʏ�/�p
�NR1pC�L*}A@�J6z�n%���U�3��������ڙ=��*a���V�ͷ����`-�?'@z�>���a�+H�C��78��ҳ^o��vW�b$y�G.��{5A�Q2�tt���sE�2֟W��c[��g
��^�d];�B-�e(���Ɓ�Ϫ���q����QɄ�]�&C�n��%��A)��� �n�?,շ�ZX4�=���Ih��;��L=p_(~�� �X�|�q"�K�s���Zt�Q�DN��q��eB�4�Z������+�:V/��b��E˘tz��7�|��}+�Ճ|��3�)���[z^.Y)_��>=�f����5��s�5�1g,�ٷ��n_����K�uGŽ[�Д��󃑗�O�1_��:�Eo�8�yn�5ǾJ�2|r\���k+�J�m�Ι�f�Z���7A�t��ٍ[��=���X��@�'�G��	��>[��|AQ��j[6�3B�N�����O@ٜE���s��]�*�L���H�}_-\�~Ř�;J�}l��k�S��5�/�V..�4�ƅy��w�<���P0t�:~]��{>�����|��X"S�Fx5�c\"4�,0A��ұ~��}3��ޖ�屖��P�4��7yf�j���v�M`�������;}��
{��~�v}A_��w�_P_�%��r6����W�G+|�����93��~ɺ��h�E:��Z|j�P��x���H^��M�u�����֐��Fm]=K�����P�cS�^s@�/���	|�"���6�J����'��`[U��K]n&�,�,4"���&�/a�q��y	1Q�Sw��p1���"]�X�"�8P!��R m<��jAVշ���{��愜�v�&�1���$F�:Z�E�VZݬXY�22^�OIκ_�����X1:���޽��4ߟ>��(�s�1Ge߬�%]p3#i}��{��]K���a����퍭�1��/��Z�3#"�����Ϡ���������}�
�~眧S-]'��������F���ā`J��s��Ԝ���gU�k�⚞� ���|�%bPo�kDWn�y�-�D�vz��`�o�;v9�����p+ָ��a��` ��7n��_���:Cd�߳��l��`!0r�d�������`]��(qfSm]	��M4���$��ʌ\Iٍ�MR�����ΞV���)^����� ��F"��cfa_�W��j�{�ӏ���O~��M~r��D��i��smDb7L����m�k"sV���ߋc-�����[1�5׌���p�-�*AFI�r�SI�ɏ�t�����\���X�;���z�Y�Z��Ԇ��i�d��l�ŋ�����#�kl?.q�&0H���$s=�q�a��L�#�f�tZ��>fH�X�]�\�˦�H]<���|��Vޥ�d�W_S2)I������E�i��<�)!�	�xg�x�G��<Y�g�h9*�m.1�ϝ���m��iP_�W���6�)/������إ&�2��͊p#��v��\T��Vv��]V�5�u� ��]V��˝jM�|��i ��Q���
���A�7�F�/��O\�7�'���V��ˏ��y�{b�o!�S=��&燠�o��7����)�Q�/�1r��FF0x'�����l��TPo)�`QiS�ϫ����e"�@UBH�S&*k���0ؖ��w��B�]\?o�z�d��i�	m�oM�zo�P��[�
]m������~{hG]�b7PH��~����jv!X�H~���l��\�hL�C$��yG�Ƙ��K�ފƑ6���ݨ��N����$�~a��}��O}f����E+���5� �-VD�RWi��3�
���z{�9��h��ڹ
�o���.?'d��hkP��^����	��D.֩-ƣ�8-��\��ɹ��h����� ����hy�K�4��ďӯl����C�(�q����O�&�QH�d]�ks���{�^�'��^6�%F�i��Q(Na�Ӽ,#�a��ws��Qꉔ	��A�~�M��Ġ_k	^e�K�!R�_G�X��N�������Z���K�N���L@���޶��/|�P�̑X��(C412�����0�����q�~µ�i�A�faL{���� ��cQ<rDƮ�����[���[����=V.�ča���Ț ���J����������Ƹ��F|��-S�#u����;�u�Mj��<;���	ho���0'7u���>P����8[��M���O'E7f��X61�X��I���M�ť����|e�鑬�R��ں��jL��ǁ{�XO��5fQ�;*��%W��MC� e�m\�{{�-�} �W9��">�.qK�4��a��������I���j�w��=^����m�/�Y�	V?��S����bQ����sl��*���Sh���m��1�� ��Yl�?�Zg ����'@ؿ/<�(���p��{L�[�1�E�Z;�Q8�)�]��D�q f��V�^�<�U�D� �\G=�t*���)���0�Pe
?��P��ˁ2�1"р�"�,���ȖDE_$jؙt����<�Y����8�~��#]8"/����C����9��͕0��/���!�ض0zq,��5�6w�`X(��rR�wi��-������;�z9�_ǡa�7�AY��')�f[��|ڮ��k���?���/^�p����r�r�o����?���}�++�I�XXZ>HH��ݜM�l����o�l�=\�*�d����%����]2N���[�5���̞$5���C\`�FpFk�(�b��R*]�t1�GΪ��-H�\x������c�4G��j8r�(����IB|0��w��E*=E$1OԲ��tI�>�I����.����_�8���~�Gtx��6���@��KUVa}��	��C�w+z���f����mZ���j��.�"sB�`��Ѣ�f��&����d��7#.�щ�8O�s���ޏ��y7����ر}4^��8����f�C�t0Q�;��4x9<���?x�>�s�O��6�m���Az:�y�x�y���wç^x�dn�h����;cYo�(嶇��^���Fh#(��,Y�jՑJդ���:U=9�TLXb	�QCD��ԈL���{�lc����S<�<� :�׍���L|`�w�>22�4�ga~3�#imb��c����p ������d=)5ۡc) �*2�E�7�9n��^��{�`f��P\`���G��W�����v�C$-]���4�?z�����"�#��Q*>������Da��DS�}�F��w�j}���BPk����B�Jd���+�V��{�e~�� 
4�F2�T�����~Tӊ;H��cp+�tw�6�-Xo�&!\��ow�pۜ�2��n1�<z�N~�3ڒI�6<��e0Ui���m�K��Y޼��t�E���[��tv��4��?�$�(��!<{�\�R�t�h����A�_��g���K_����(�?�YpgX��d"�y���c}������E�)���I�Q�*3��j�{�1��~�����ޙ�a�A>���3�<~�ګ�'���Sa�e[�3�aoC:o�{���a���FN�Fl�(�N�� R�7�I��FaZR����	F
ﳛ��&2{�$�#zW7�T��?���g����P������#z�x�����;�T�u�9��u���)6˕b��HY���3��I���Wq�&��	��ut}���x��ΨB|�}��;��\�"Ѱ��W�a܇�ww;?���0�pa׍��Øvl�J������$y�kX�������S��b�u�)� �l�xc@�����eu�����_�z��q��Er�6�}(�b��t5op�[��nJ��;u�NSs[[S�<�"�mnšV��鳡���G?y�ݘ�Y�@w�,
D�M��9��1x���BJ��`/�^
&#q������!Yq�QH+x�kh�[<�'��tpMp/��>L��~�0K.�f������?A��O2O
�>��H>)�]���p�Q��m�Z���zژBw�Y��pVמq������$3����2s{����0s�d��T�)`��΅�S�����p���%P�-�G����NZ���g #U�H�09����D�Ů�Ţ�.��B��v����ǳg���UzKʔ��0'd,l��{�\9t#m7�ΜS0��T���M�G�v����s__�۠Ge�D{���ŵFX��p�(���>K�-�M�s��J�c(���O����={���9����ZW��b��R$
�#QbّoG�2��	����:�K0��Q�@���׶�`,0�I��|�*k�e��!��1�-%{.�P���F	�����v�cG��~�d�Ma����VB�$e4�S�e_�H_��C3��v�M`6�o��	0�G;���N(Z�4.V�h��B�m�a���s�:���P�֦ul��"��C_a>|��ݡs�j��2������б�~�Rm��$��7�w�TsX���'���C��#P�<BρP��6Z������r+�p��[P�ǆ��,��o�h���u���{�gz=	$A>1��F�f����.ݝ�*�I�!q��%�z�v2`��\H*�f�����"�Ab�*�<�`dz�ƴ�y:,��w1����q�?�ހw�~<K;M��1��2S��_%x�����hD�n}�ǯ���?�GPFP2�Ѕ�w�Y��}���+(�u�bo���6o�ݱ�a�sѓlb�E%E9%35�R��᝛�e��2�Y���=b�r'59@��|p.�������o������6��2(}mBW���J�d������܅��,��k`�z�v�{���+_��w%ܥ蠃|�s�}2�-_c~z�o`�]�ەnc�e�G����eș�U�[�k�����R�O�wƽ����i���e�!�(!���X$��L��Q����$�*��Me���v�l�.{0~?[��@Ý�˦�KHꗸ��к��-"{�����$��R�&����Db��D�S�#"K[=�l�T�q�CgU��I��*У3λ�o3��{v�=L4�_�L�^���Z89̌�]F�/pO;�xC�qLr�اs�[(nȘ���e��>9ȼ׋ �y��e$���i����5��M"M��`	̭.�Q�:���Y����h�[��vEx��B+^�
�w�~.����3�u7��e�k�>H(�2IY����At��H'��pm��q����N�����L�u���1�I��סn�8�DľсPX��"�ӳ7�w����^XQ���^�t�%����0 %�]�$��m�ݏ���k���D
���?��Moq(��-']�^+d���������1}���0�5���'a��G�0�Y?F���uQ�Ï<�Q��C&���If���gyX��'��C�hܸ�5�\t�����d�
������#����D<!������mf�l�|+�Ve���͙hs.)�!Da���Ъ�� +�m'Y�j�s�ys�I��8��+B[*D���+UH�J�>h`T�*L#����MiXT�.��\˯����*��6�R��H�dF#3d�=&�����Kwc��Ņ�����vtİ�B��rh�;4z�s?ܽ'|�ӟ�����Yf������f㾗��x��µ[�)ؠz��ce������I)���>���|����c���;�*v�SǇ�+�}.�����O��cpy�Kk���#4N�X؈Jc�����E�5�v��)֋L��E��SGO#ER����l�`���.��I=b吽�oeW�-6�Q�0h#�Z�㏆�s$z��'>�Hx�'?FI��O=�,�)L�����(b�kc�D�H7�T�.F�F�:�M��Z�&�s��ѣ��{$�w�P�Q�Jo������&�_
7�.�����;{EE�T���U���A���_?�iς�-<h0:߇���sf���\��ۿ����ǆ��Ty�E2�z�)�+��Q6{�JG�h_��V�f�;Ņ�*(�0s!&�Qn�?6�m"�}(�f`%�������D��'T�eTS�{0xN��)��s���f>Ӣa��2�>�\�`"џQ����5��Y#�-J������(�B����g��
��Dbȴ ^1�u{R�8^8VE��ѽgD�ʚ�g�K�υ��Iɖ(R�`�b��F�N+�1�S�\`�)�&������}�H�)��K�3����+�B?ԅ���l@%s͝��1���"�`��}�(�H�1�f�7X~�<���s1Y� E�Etm�#%�ۮΡ�7�������fe�[-����R��4!z��ti�P]D�I蠡��6>�<�=@M<��h�8�|/��ģ���8��v@	%B���L�@M6.1��Y�S�A�$�q����$����-��?}��d<��4Gϸ�B���Dh�C�R�B%� ����Dt��,�/|X@Eԡ#ǢQ3�<��� ���_�z��|'�.MUj�C�@7��'=�Ǽ�a������~��oѝ,	SH���C뫿��3_�*=%�Q�}��An��A���J�zKom��$zkS=<t�8�ٍ,�ߐ�Yr%�@F��T�a��h,���
�%��F��
]�*14;ͨB,e��X񣑖�2�B��2j���b�?�s���,T�0wP��DO��ɻ��FE:G�[�	͔H@���k�O<K}7� �H&�Әh��5��vr2��{�e��*�vh��ʨE�e%�H�y'Z���;�W�z,��Q}��9��"�Q��ڸO�C��0��z�����r��̙��'��3��H;x�0���{��y;�f,�3O>#������g��}�0�&w���|�f�73��跃H��Q^ǝ��,�J�&�d8�(�1*����󮥢�k06��Ю ?-�ٖQ@ˋ$�x:�Q��((����k<�ҟ;Mn%R�3{�٧iz���_O�O��hx罷c�G:�fL��/5�����µ;�Q!s�)�=�S�R&[=�r^�.�eR`.�:��]�XhQR�@g5`�m�sW��Je�wަ�s7=P}x�
^���,3�g��* �Ҹ���E�>��\�`?@`�Cf�~���"|������� �.�"��������O�5�<
ὓw�)���T������!�8v4Fi�@�4�bc���?s:�bFv?e��(琓+�F`��^���d1��]#7��B�S'���/��0,|�ʬ|>㣡KY�;�X��j��ׅa�wT��l��UC�P�R�<��S1_q�^�a=��g���w�̩E�8q"F?�1r{���H�Gʾ���ш�e��F��U#� '� �r"���ω�~JZwb��:ڍ�v����ʨ$�oj<v�JE��98�p�d!�B�M���1|���ӿq1,Q�p���	�3Uq8Vi=��m@��ۣ��"P�e�����>����O�s�v��y���=FG(��DTz��?�i����_�HnSEu�J�N���J�Uч\/_�T�;�d5M�
�j��z���c_����/��෾~��_��8b~:�3e�aXb;�?|���
/�ЎS�B��F�d��v�S>p�@�x�k�͋0���@4���D���y��B�ƾe	���(AF�N0m�ޕ+���5B1��mX��wh�����D\	e�OUM(�M��Y�M�&�I�7Pd�9��7)ٜ����_�%�'i�aH�{�����C'���wχ����a�z6���5r��߇RZd�m7�k#�k�خ��p�e�q)6�!�2�>�t�nʛ�@������1�{�1NŮW/�����Cv:�w�퍖�6T�^_�>��2�#�����I�
��E8�~�������� �Ed���G��7'��~����1��QQ9_�P+���B�|��e�@���O|"�Ǘ��*�V����y��نsb���溨|��5�������-ȸ��+e�*�O�u��U��1)[d>��� �d�}ᙰM���s�!	Q%�OQ�繼�\s��Ң�g�J��$Ė�a����^�%�8C�y����y�����p����߀H��cp�
������:>`���VY��H�xȪz�<�����x^ �;�@!*����W�B��#��0J��'��;��7�bd j�6��*˽����R� ��(����|�ʤ�����!t��HE*�N �$&I�B�����,�E��ص���w���4��)ɦ�S���(��,�.`�6C��@��6�B؍���^�NZ�h����B:X�n	o_8��"���BJn���$U+E&�QB��[?����`�N���� ��s�~!,ap���=p_���d��ҹx�<�f�m9��V������o925v�C%�"3�_Qn�U"���z˷���}��sYR\��J$!�^����^"¼J����ߏДcu��o�f�r�R8Ŕ�x�ɭ������\\=��?��m��p\�D�~w��Y�3
��T���w\)]��~_�P�r�V_ y�i@��Z�&uH��>���U�HE�|{Z��8���-�,e�`�����6���\�����<l�_��sa���L�p���v��뙧���w����?x ��3�|.Vk)��}��HZ ߙ�D���w�6�$6L�%�U��$W�f�b	d[����b�
J�I��#�w"�}���d�`����X]�/�w��8}m>X�����3t9�rgW?�a(����O�������i���6k�Ä�w(MR��2Z!�i8��h�z��^�I�V�q��<�x�h*���B+^���`�[����+>�k�9�K���PG���$q��(P��.�7m�#�^�cl�V_/���;�gV���0"�$�m,�W��Z�����:3��:���w�
��9�Y�$����,Q�P�ȱ����&�M�3H���"��(a��:�on�&�X�s>���2�Jk�d��ΰ�e�=Οzŏ�Fs�aD�QПf>��N�\V�0#�[�XM��(E����b�`��7a�����GY@�W�
T��y�^�!'%o��Jdҏ�7rj� ��_嬢3z���H�+_�JL|�f���*@��U��ynݺ�o��C��J]�*�Y�	8qq}m�&���u\���w'P��ё��޻�(�D���8C���"���{g��j!G�b8��1�cZ�mu�Q	��H�SP�Ĩ��5���R�q`��EX�e�Ab��n�	7gW�ʻ;�
7��6��:�%��H_�B����y��kK�[:�q�{�>���ȗA���$���}�� �Q��G��o��҅�w�����mP��E�y>o�@(��	��
?�ᷛ��'<��~��u�z��s'�yc�����y�����������~뛓|�����9�v��VBQ�v��_�瑩�,�`��,�	���-\c��^�8���OL�u%��.�����;6�u�.��P�=�r�*���i� 'l%/�<xx7Y�(y�U��؄.��:���������/|��o0saWG�^�t�������}tϱ0;u^���$%�o��V��9~<���k�c�9v�A���z-|�O�a>�P$(�&G����Xk���9�̴���꭛���~0J7��n����Ȣ����k�`����w7\�)�� �L/1Y�uh�.��e�җóO=��e�^+'�L���Gq
sh4�<;G�-�X�θ��{{��;�UGx�v��Ra��;S�(Pؤ��i��z����o+��~�~ B8}ˍh��cǩ�`.B���6!ni��<�б/��Qj������o�c9r�HV���o��v��W�j��څ��ڍ,n�Cc��S�����23!�/���:*�j�tϪ����Kk��6Ո��<�,��q���a�����m���]b�OB��;?�����>8��M;�eD�1��m����v�j���]�A�Zta�)�!Qv��A)ʹ����<�O���;�g�}<ݪ�#�(�2���bՀ4�o��(��.7������җ��Ƽ�*�Q��wn��pW��s�?��Omp���&�������ױ�������ȕ�n��{�x�Q%R�1a���g`�^��$8��2z����R;y�}�����S�Ė�M򀭆[����lŀ��P�Λ#Gq���,F1�4PvR��87��ӟ�����p�� �J���6�~�(�����\���cxć�6I�}@hSx�C@[ur�wn�q�����o�o�:���ù��Ue3c\+�~*���_�e�������A871:�;&�^f�<J��BĲ�q�P5HR,���{=&�Uv�����p��J>�����C�u�	����d^'�OS4���3�%��7��d��20C�P����O�o�z�˰��7�K��X�֌ ���k��4�M�����oKL�<4<��?=s�dއ�QSYc���l��J��7ߌ	q���HɄ���H��۸�w�رh�w�}���p���s�h�|.VSyx�5PǏ=����j�Np��9$����8��=d��ӧR���e�a�9�'{P��鉎f)��	>.S���� 2+p�=�p�֏~L! �i�h�|�R�̋/��]��-����󉧞'O��ƀ������Hl����xp&/�8T��
n��z��2��&��x����]ݨN��oL��:�rK�ֶ�����]���8���޹���^մ��9�b���V��ɰ��A��jkjne�R�*� ���c'����7��j�P�;ZFyL��P�p�HTj*t�%e~��Ujq��M ��Y�.p�*�e%)<�(P��I�`h�ƞ�����m<��tz������;��K4Lz�*!���*�I��6s��<�LT�Μ�d�+(�Y�S	�� �<Y4�Mr1M|���_!IN��쓏?��I��d�s�j��b9s�e�=x�$�;�gU
s�% :�tt=}�s/Q-��=`��$����2��/}9F@��x�8����$�O��-���U=k��U�M��&T���|�]�Y^"/A�
*���q������^���R��"��
�iМ�y��DA�4F������p�Έ�iT��*��}�Q�zm\N��k�A�hk<n�C����*�ow|f����0�*�}����v�F4;����4���������ڃb+G��s w�u�&G��8�w��I1�,��
��xjn��c2eR�����Ķ��g)���ƻDB�ר��W_.e=���2�Vƅ�����ؗ���N�EK�Ji�d;T� �{�?��s�]'Q�~�Q�������27ba3�!۬��EmtWEo&ٛ�K-m�.׷k�ރ}�]�^�P55�\+5UfG�Ə��ڽ��������������j����-�EK�-C�#H�FEQ�¡�R��
�\ß"�k�o��|PMT�=Q��S�������顃����7o�7�x3N�ӻ�д�QP!8�hj�X'�{��d?�p�x�vT�	�νa��4�-�B������0��N�e������q�Ng�rAz�T���4��I�}�2lmf5�Β�$����萩6���yZQj�y����W���z��pp?���3��ᇯ�����[aFț1q���}.*jYs{���%���5?Q�����d~޿0,g�����H�h2?5/�͚���|~W��=��@N��9�*I�lTo�\��J8��nRn�Ca�J��@��gSa�]Ow_�o�و�cW�߀�|�l+�4*:/��B��U�>�hT�F&F�q�͂	!��z(nW������Oo��/��/�W_�q����.�K����^1����hMgƱ�Q>QF�͌��6kh,�󉕺rtEZy��6�=�LY�=6U�Эn�K�:��.`�:0*��n�r�8	��T�Yv���ȭ�kl��g�" �vCk��U�{ǹ.���3ɬ�*���H �1�����k����z����ɉ�X��z���hĆ�Z�{�b�����t˝��~��5��y��ޯ���(�M�O#v̞�`�u���F81�%�"���������E81�Nl�ƹ�0[x�b�B\$���0�� �q��t
o�*
�Ev{��Q�b/]���T�:SDTT*���K���K|�M3��P�6�$>��3w�wȧEվ�a�C��UC]�`�NJ�kP����|g����?����C2����Z&+.���$���;B+4�Ҫ?|�ʜ��PD=�|�h�Zp$��SE��
�5��ɶ�0� ���6Q�VR��Flm���*�l�"$j$�r�z�y����3��ǻ����2/��\􄇇�ޮ�w�}7#%KiU���2�T��e����կ~5|�{ߋ���X֪̦g���o��#��1��5���i=<�D�w�{+'��pe%k5H09�N�k�j�"��^�¤�o��oPtq&������s&��o�V�}ԟ�|�qx�e���P^���P��c�.\����~V(
��@�RٷR �3�83�/�(�`Ni�{��ql��'������2���l$/e�YU����<�i��e	$��>��5��1+�ר�F���5����k�Q*2Eu��@�Rƪ��ػE� ���f�=x�K�P6����&�#��M�>��#`��b	msKT�=0�>P�ɱ#�c�[Ý��.��w�9Y 	�Cw�>�n<Q��nn50>㑺�����n��TG�W�.���3�Y����H�<�n�<��-����y'r<� �\b8�=GHbwEMQ��9#/�cy�d:܁a<K�v�uvG�P��)���\w��<��Z	�	Hi�|	�`4bz���#�:��+��",��	+�z4Z;�]߱�#���^|t���ϓ�s�H
�c#?�,�Ԧ�>v0�X�I�?��x*d���G���]���X�\~��Ź�#܏Ǘ[�ch -����SD'ca?%�$�K�C���~���!/I�B�7����ĲQ����'?���L���9�n�o��96H�l�]ҵPRٍ5�ҶH=bR�1�0���8���c���~����F�?G��V���[a8�%z;:q4����f�y�nz��%��z��wbd������o�1��-׸x�sR�}�{WO��
����
e�2��;PY�6k���a�bi�E�^ޞc�2�-y�}z���H��f�B)]V��0&<OK+����s/}&ŀ؅\����H�u27Ş�#guhLl�;�W'��P�@�pT�{���ǣU	���@�<	ǣr7�1!jE�A�����(����RnS�|	�Mx��U����2q~�(G�������T��J�;}>BN5��-��~�9��eiUl�%Y���~�`/���Ɔ�X>��~�/̑�='�r+�g��١Ǖ0��#�h����������?��?�z/|������}�닼3c�qQ���3����Rx�9n���*�$:�&�)�Ȓ�DR���s��&+�m�ǡ\<n�+�k	�Ǭ"��������z�+͌.5zn���+٠T#�b �:f<Qʖ�=�5<���b��<Ш��%L����0��sχ`�����[�&"j!��P?��cp�A�ñA)��8}�g�c�#�S��/�����%�����ޒ̝$��y���7�R1BN�և��|���T�2�TW����vud��*vǓ.oZ�[?y�r��=�4T#�U��0v�=nGw��<0�^r Cx�4
�"�j#�|9&��(����$%����C�oͅ*�������n������@��/PK���Ku&�-b���;��7.���O��?����r��gO�nr ��;�Dޥ�	%Ƭ��T�ݽ6�Y�b�,e�1"�$H�QO�PZ��j�ڑ�)��j�_3�`5���u��0��dy=:�ʦ���ZʪQ���IYl�*�&�Ռ�t�-%�рj ��&#1�;%��R#��;Ö����V�����&�i�;��@%~�̳�NG��W�M��.*�H��:�WZV"�'#����O?�!��x��s���V�0�UO*�q��"��2�=3]�gc9o's�U��me��$�WE:GΩ:|����^���޺��b�]�lrM{?��P&Vj�12�(x�]�۷�ؙh[CV�$�~h���Li4�F$ �e}��grq9�o	�/�_K�G�7�:�A3����Y��>���Ar_��uB��1���P�Q匡�(����}����FK&��*���S~�5�������<`-xU}&�}�|ȯ1'|[^'<�E�6�s�L�)���iࠎ0L4���:�D�G��?����� �?I��A�P4Z�>k�b�^;�k%�T�2�(��O��	:��)�Z��8��&r��1o%?�ѸI��v�]�#��݌9�2S��((�f���ǎ�;�`��?y+<��O2yod�(��x+y�Y�po�i�ۗoτ�C�B�(�"��'�Q��v���8_����?����|���>r"z�vA���N�YE���[mG��4�n"� >�#ϡ!e�W��F$���7�G#���M�=f�;��Мiy�^��>�b����M��<�V[گ!,d�@#�g�J��K\h��0��ݟǧ���hC\�g�&���L����t���mx��s5��z�,����È�m�h<,�p[FR���n���w�8 g�]��GyP�����y���s?�
d,�zu�p�>��*�'��?��?��l3�.$��a�N�9���7�k�u��2�,���3ܦ���He\Rf��)�U=8Y��[����>����U��_*����ˇ��ʸ�VSν������pM�`o� ��f1,S@U���kt�-���+�ZVE�ܞ�CcPd�y����A�X��p�~<�F؇b�2J(b?j/�KQ�>p�&��*��D<0O3�E
��б2��B�_�[������?��p��=�G��%���{���wi�z~�U�� �.�#K0e}��ȅ�C"z8�*�y0p���
���ñk]�CŴ���)�/fZ�o���9�j�@e��q�<�����"��E�k@4!���#����N���T�A�c�a���F�}��U�BMvsk@\�{��y)h\T���^z)�F�qn�5?�r�{t���@éQQ���ГI�J��1�}�1s]��u<>��Ir��5tFùq�Py�ޓ9{Tܼ��^1U����\�\��l?������(��s�����'����/FUϓH7�?B�*|��E���0��C(4����z H���~7��)1ۙ0 ������2��Jm}�T*�>�.3MI��#{����Zhl���!=|4z쉰���%�N��)��u�Bfa:i�UvtW(���,��\�N�i�߄x'������~�O�oBwAő����=���3����1 �"TAB��dl{ȣAeс��F�ߦ�7��������^x��D��[ƞ.�;�i�$i<f02�r&Q�Ti%�T�,sx�Ѥ���p���J,hF��]ԋ����%�0���YN��ɉz���a4��'Lb��N�;/ý�s*�ι�s%�I�����h�2��o~��0�c7��R��<56ߖGEId�T���<�Q�Y�����}�;߉�b�# ��\�=�V�Cc.c��FG��}���)��ф뙻�0xoi4<n[9�����~ܧ2͍�J�s��ݗ���#�Gq@.K+��m�����/gtl��w�y���H���+P��2x��d�έH�)�X��������L�h�65�N�܉p8��T�By�lZ?��~\�np� �	�$����֫�Cq���@�Di+�o� �^���x�gHP?v�=�7-�7Q'�)�x���v��������=��
�cd��P!")�2���_�`n`�ʤ��,h7��Id����V�ʙ����c���)=�us
(��ԡMW!���W�Μ`��ѰF��w^}/�7�����������.^�|��1���mLB���4��t�U`[�k�](��s��QSq���D��c�.y!�8Ir�
�+oG��wy>��T����=��S�o,1e�9�S:$�$�aՒ�M�v���/=2��j(�3�Q�	�$��}�{��Wy� D�)���ܜ���=?_6���E���x����Ѝ0�
Uc��]��}h�~�ĨC��h�ܗF�c�{�Q�砼�t�M�v��}m�e3eHnt����h�=1y `���>&Ɂ{��H�ͮ6�6sm6�`���"5��2GY�͇N�}*��pF{�#ً۸���$�rJ����l��mO�3��)h��
Sx�����#�
���������{,�5R�a��g",����_!�H5{d�-��*U,�.\�#�Y(W��V���d��d�0�K5z=�����0P�4
�����݇H���*�[�`�]@\]P��}=�ݥ�F��a o޹Nc�OCF�6���I Y�\&B�;�p�A���R��9c�H����������w�~/��PF��	o�q*U_�+�á[�\5 *u��U$�K
���PBGULK�w�W:�UQ���ͣ�i^+�b���E �^��\c�9*q����k��S)��f?��0��xn�eT�z���<�1B�\t rZ����^~NXń�p�RW�O�����)����	v��5�����x.�G���ZߊFw�B�e&<F��r�&���]��6Sf���46P���W+�����D�CG��ѷ����Pa�˕[S�O�f)Y�s|� ��o����up��16�ۂ�F�G�"w�c©�CG���	�z���E7�Rh��J�+�A���ټt�]�@��}��y�n�eY��Z)@�19ǜ�Y�R
���Ka�ϫ$�'�À�.�ؔe��-8��*<�l{��N73H|��"��PP�5Pv+x�z�W�Y�H�:M���Π<,�5���iρʩ+�"3�����<�����y�+@c�8�	�u"�E �5��2}'E�'��T��lg�sm�_`*#�[$bW�t�37{�ߤ�Ű��!�j���f�#}�͸�B5�91��|,�Y%��<��a��<䏺���\��%m<ё�V#��?	�3 K�Nz�ۍ, ��=����L�w�N|��Z�х/=�<∓�P����z���w�̅�����o<O#;�ͫh,���U#�65VDNY�Ap�FHc'�Gh����ı� eE\y��~��|g_��N���y
�50"R�oK���9��rj�E�^
4�r_ˡ�l�*�Y���\���1��v��`�Iz=(	$��$y�Y[]�#�Й{ĖH.��}����<Ѯf�M+�TzS>�6�!�kŻ+��W�n~�v�>��>��^x�x�3�;���=��0�L���]tQ��$��Y���q(�8��U"�B���Ӝ'/���Y-�
��,��(�/K(p�ׇɵ�YǨ�ڐ�c|5�o0�ɜ�:���`�4�9��v�2��6r1�K��R.�����'�}�/�+���f��o c	1�Pc!�ff%ҥlD%�b���>od�i�w0o���Z%�5��܊��a�{���#W��a�*�L�g�^�^Rii$�BV42Sn�o�`NCn���TQ{�F*\��W^��~�hE���&�����U��o��{CC��JʈA��}��0R�K]e����}h ܖ���ʪ�v��ͼ������9�y���y,yT�Gm�0a�����$�H#�AYs�|��c�ZF���G��0���$�� '�c���Z߄MXH.�l�����'r�e���	M����cx�7�n��2
&�qUx��*)���
!k�ڡ�����:]�*����G����k������cᩣ{�޾ְ��5�Vg���D�������L��,S�ڛ�X���vŋm�s/��0��k��G�.�Oe�]�۰Od.�&�L�i$E;0}0�6;[lZ�sDR�A����.�a�|�VXQ��,��!�D18�jY�p�:y��6 \KW<����0�Q����ԕiC�s3$Tq�k��GU~���~�!�{��<���('	��1��a���Q��b4!�79��ܶ��B�̗����3��G�s�Q~�ؘ�r�zپݧ�i�T�OV�����^'�R`g}?��M>P�a�ܽߌHtP��0�.�����O��-e�Ar?�#�>昲ʲlG��wTn�������Y^�x�qLt:`�4+\���A��J��{��\�(N��9�F�b��Zi�������i�d��(��	RDT^�o]H &
�P�#F����&�v�����x��4M9�o~��b�	���7�g>�$}����]P�Ӹ��>��c�/=>��'�D���ZX��n���=m%�d'�h��/���̾n�:*|��A� �Wuo�����yw쪵����_ ��w�3�"o)�j
&Ze$��9~9�J���\%|�&�� �`av.~�;���[7�B�Bi1��JF����k5�#}� e@���*��bʫS	��~i]PJ����@�l�@�8�ԽI�<���4T*,��e[12�X�.+��uz�F+��X	x�*t�hU��OY�Y�>���H	��Wi����k��k�r�*i��8�$+Ԥ1�พK%��VF�R�Yw]?g,p{:)�<r��w�s����~��xnnC�,/��i��'C�������J��Mrl��s��C���?)�w	;��2��Jt��?��Q�[����Н����1�X�0Ѩ��l!Kλ4���~q%�sk����@&ov� U���x`{��fP8��xX3(��7�"ʨ��omuvy���;xX��m�f>xyx���xغY���R�TuyʘQ`�u�q�އyfvO^�]~���WI�¬{ �\g�^�^��ӧ>�nĐ�3�Go2���ՙ�m3�&\Q�?���d5r���޾����X�uF��u��3�Ь6����U�����N����NM΢F�<J����L<}�\�,g����r�$з��$��2��l��Ý��Q��n`�|�s�
Ka-��r�Sa�<3)<����24NL�Ô����#wq|�Ŭ :��U��\q��Ϡ�p�lo������竁ț��(DJ�XR�Ò�WY��x^=t�߄�5o�S�OP	f����Ḿ��#�>zgT��#T���ލ�Q��g�L�sQIkH4*���&���4&��FJ�^vh6T��Q��p��Q���=��уJ�(�R[�������<����4(�w*n�U�Q���q�h�<��%�3���Q��Dlg�O�_(o��d�U�����p�����!����7��g��ʨ�'o�4;��1hh.]�|]� ���}m�N��zPH�I�|�G�����������a���6Ơ��h�pCU4�M��fYCԴ\�l�o��}�u�e�(�VB��.��^�A(��m5�X����˕�_���3H�f���?�;;[(4�Y=��H'������x�y�YU���r@�jx��M���#ǥ�A'��O^��HC]m�⥳4G�����d[���.��ahЁ�P:ܺ�T��A���Ha�L"^����95
�h�ģ%�E�� ԓ~{��E���`�-��`Ԩxr�h$$�.�T��$&�3ꀆ�Q��J<��>J���Ѐ���S(��0%.Δn�AI����KnbZ��}� ����bk�8�6ٌs2l3��{#��xd��Y�`n8�.��׳VY���������Z,��9�$T;v"z��㭱Z͆�<O���Qp2�ЏP�Г���t9����k_�Z�P�j(�)�th6hi,Vm	oi�ݎ�(��L�������Ӱ
w�}���,��������Cc$��a5��z�^�'r�j���{����2��8�iZF�D�.k�����VJ���B拳�51�R��P�B���iفz-~h㚴�7+[�]ۆKkk��A������mc����ފw���Ԏ7_�+�@e�QDn򦈗�w�Y2�bE���wn�R�Y�nb�R�
E#S�LևJ�#�
��`��A�e��ڍ��Joo�4���:�oU8��IJ0�[C����íw>BRY�O2���R�'�/0�����Ξ;�I�ϡ O�q��l�^r�=�t�l�����Fy��]7��KG��Y�>��B�� �p��7n^a�&C�����X"aN�9
���5�l����.:�-�UqA�}��y�j�4��l�;�md��3��j�(���c������B!X�:�����������l�v3�C�������$yz�TE�b�c�h�,��w#$A���{;�-+ͥcr�G�3��bBw�_�qX�$���E!����h��v�0�
���m���ChD�w���J4�]�`�A8���[����� T�q�W���4<���ϻ�݆�׀DFl^r+�����T��ԅ��ba.�s&�5>/���8��]�-�ч9��8�+ϼ���u82 =k����H�)���R���>��-���}�= \��9����u��2�Փr��%Á(�?�N������C������u��D�r��4��Q��A,�o��`�C(~��B7T�n�q��.N4e8���f���T1ba���������`�����܈�V(4߸q�q�L����,��`����ڱ�-��Q	�iN���>�JdP�a!)�V
x}�TI��2}*���M���Q$�4�	_��3P���"+̓hb+����.(KJl�����'!?d�)�ޅ[j�dyc��'���EJ�f<���:0I�ޡ1��I������@�H��� t�]e��v�NH%.Ɖ$)�pV��
e�\�Q�=��F�|��$�ۚKК���!���b��N��:�e�B�E΄�y��YU�=[���;P��"�=�Y�ʠ{+�\Ʒ��D"����!&j4��F#�$$t��ur3w��Nc`����K1�p�*q�&_rB�S���={���w����8iPr+�&��s\吏Pҳ�>��у�d�����n���w�#�In�/a(+�r��\��n�όX,#�`���8��vc`ލ���0_�sϣ�����;���-�Q���,����1r����t�U(�h�9ǽ����aﱣ��pi���0��r��\�7�{M*�b�Oa������AX�d8�bw������L.X<�8E���������4�����K�͕�Ɓe�(&�C�p����Z��@���J	/�[����7y�n����x����ċm��|ZZm<�hĪ䴆�����*i��os!�"e�ehE�Yw��+���{���x����s᝷N�٥ס �յ��H�&�����"���`H։\�g��Jґʕ�%�#�H�Q � �2�餪��H�ԙsa��=a���l���r1Mvc3K�@Ua��Hñ-EH{� ��w�$=F���Ԥə����@O��!Q뫋q����}IS��Xa�����ьIn��2Z�T>%M���x����P��̿�6��������j6�+�T؟x��XY�qJ�E%}���W�Y�m
s��Գl�=&a0{�z�ma8�y��FHů�6���V�]�SmI>�K�29�z����bԠ����t�g�7�o�7��߈�%��ʗ�>����xn.����N�4ꊝ�8y_Ln8�j��gF9��T��!�W�-5k4�?E]Cf�7���j�`�\�۶��Q*�٤yv9�a2�m$��"�ѱ]f�rb�{�|������~��i��Y�q��O�l����j:D�z�V[%8�A�	��O�J�Qe29���W���p���w���]4܍�Є����V�ȅ�
 ~%*gf��Z{�J�P��b���+9D3�0���L��40A�z<&�Bo4�����ڈ�s>8}�f]��3�m���^�B&����BF\��r[g��L"�A���Q��Z�'��ŀ~�Q�
,��D+te[�[��6��v,�b�+�cG�l6"U��>������6�u"����(*��01�|��*�|�.+D94L|a*O=�2r�Q�!s�?�d��J�0<bz�W�]����U�-O8�Ǒ�M��J4��� �����G�5��f�W#�$�e�DX�>���I-/;Vٻ{>���*�c�`D�[g�|\����خ%�0�r[����c���e��4�^��#��:�K�q$A�e�c���q�{4R�y|+:T��^*�۩:Ġ� ���H������&��8�@�U��Th� ���nj��Y^��7j�a����)� ������Ю�̈́;L�y�p7���nޮ�uJh/.L�M�2P�*3�@1��?�q���zmu>luþG����#1\Ә	����N�8�O�Lww���$�1�����Z̋���1ֵ+�n�*�M��.��1ob��ʤ���� �!�CQu0n����	(	�0��:���k$�c�:��AT�	$QCYlI��n��F+F�ϲu�� �ki��b`(�&J�Xl�чbc�N��m�
��]�ȉ}:T���<�|:
�
|Z�t�#�m�R�}9����9�Ü�o�SՋ3��#�|@�X.�!��|vhԫ���v7#��m�K�iF�J5�����չF�o]	�Ξ��r��/%�J��^�ϺP9i`,�ի���.�γs4eN�bR�!&�1��y(����}x\F"�<T�*��V���èh5j.c>#/�5�1
�{��|��M�36>��C��QC����2絼2�wS�@4�-f����xܧ��-��p¾���_�sOu�F������7��0fѶ��:	VY��<4�9ߏ�,�x������g�#��I�!p�1Fח�B��mH�#�;%�͝=���6!iz=(	$��$yۡ����=-˫�d��&+�,'��C�%g�`��jOC�ϐ�ev��#]g£0�8����Sgß|�����4�	��c���UǙ˷�����(����.�}6b2q��
�����ӳ>~�L��,���o߼a��������#9-�
��|C&��w�$���*���QoUYw��\6O�P.�1���&g{5�a�{��g�qouԽ�y�a�qon#�!ɿ�x�(&+�퉞�J����
�X�1Z�����b*��r����)���{,'�7�@�lT��-��t9�{�]��(@��~�0�f�"A�����ܖ�분t��9;�2t;�C�c��Aјyޮ�ClVy]ݧ���<O�����~��j=�/��]�}�;�������"%�ZhO[�f��=�6�������e��"�,h�-�2�^H�p< A��f��L8}-!�8q~�p<@OR�2���VÙ�+��(����W7x�0,�C&�~��6���k�
���4��?���������o���^�.�	
P�w�I�*�,6�b
[�h
H�ġ#�.�%z�{�ÁD�Q'�v)��)�������V������>���em�S�(>LH�o��5�Y[�'V��}�7�x��J"o&T�IM��P���*��r�V�pEݛ�����D43,����kx��R�S,%���h ��J$��w���_��U���	I������Ө�-�:���V��6�M%�rV��G(I��=��+��6In�щy%��|�S���4��]40n/o��xN&�U�.�~��rJ���(s���2��cV��r�K�s�C���?e	We��a�d�a9s}c5��Ę�����{yDc����)����~�Ѵ��J �����h���[.(k��h���j��q�X�=D;�T�=)�~�����C�����L�ٷ?<��2�;�i�����ù�wÙ�Ӕۖ�F��Er'|���]#�۽�~5�������r�����.�K��-@A*��@�p��U�*?��^�gN��y�T������JLzta�H��9�ë$64�Ze�JAE�UN�$�Jz[?�Qx,� �2Տ��,��G���Ai������������7�Y���G��7����(�v�|~���� �>�d�JO�k���ʯĈ�s�,�D���jx����N8)W�Fn_�nn����)@<V��Q^+�jD��h�L0����nt�㱺��L���l�̜N>APc�1�~���>g��#����o����
�8�/���%w4Hʻ
�}�S���τ��k�01R��P苾��7����@�<��!�����Xз��UF@FBD��>�W脵;Z��"Z#Ґ�Oe"�tC�'�,�ۉ>�n|���|��d�p�v�z���0��e�����>�e	j�!7���no*�fn���V}��9���M�5�����*�󨍉&n@5�g����^�R���{�e�)�4� 79[i�ċ��"K��^i���LF7*s��+#_NX���ۉ\�drÑa�[����9�)�#ˡ�<����;�U���
N�.�޹��ޗ==z���
�DwN�a���r6�!TA�?�5���6��s9_y�\+��~������Ȉ�ݶhP�B��Q���#:#���<?����=���^��q��Y���<�̨?�F�!��u�*3x2��2Ü��� �n{�}&� ��LC���7z5'b����ǫL�"LN1�Hv����TU� ���n���mƚ=MЇ�'��n��J6#���dT�z�+˙7���a�s,,��e���X���d�Ӊ�}1|�w���T`���j��JZ`gM�R���C$rsP���� �E` �%�z�����
�q�:�!v���/Eá���vQ��m�2���C��[�cPx�m�3���;!UTp�K��1���m�����k��΂�T��o�ӲNr����L�� ��Uڱ�+�r��i�b��5���Ͽ�B��Tw��zF���9�c�fn��Ͻ�X�c�q�Ʀ\�l���|Ļ�mDE��.���.R�Z뫏I�rSid=~�eft����!�w�n����}��Y�g�ׯ��w��9չ�30"sn3'D��>��O��}���@hU�Q&�BC�_��èC�?�l?�[1�����C��#7:y~*7yinfH��ݠD�l[d=�"��M��l��F���AO�ۑ<�6��&�	\�|�~�a��T�������W�2�a��zPHǃ��}l�^`������P�(,a;��v�-7����k����QBV�H���Ï�\ѹ�C9˃�|�Th�j�x(Ҋ������Q�����{����_�����&y����G��DU�a��$��/Rd�<ʔ��
J}+T!w�C�T�*�8>�6w�*T�x����1�ѻ�I���w�-�Qa*�{�"%��0�JVl���K�"ͽ�{s^*�}�'|or�����/�'o�+L�GT�i���5�0$���m~FxGe�l�37rTQk,ɵ�)g��h\T�##�э��{ÿs��~� |���ay���8ʖmh|4j��b�����6��r*��^o�Gc���)��F>��}e	���sy%7�1�"�ٰ���S��:-�d5u��PI�,��q,�Nт%�뇑"��M����~~�d8�0�M��c�Ɣ�O���D��UQ�sx؋tB��Tv��%�Y�`�s�ÈK����s�������3��������u���+�ay���w�� )j��l��?�H3_�Ik�eV:�\�{>E��E�౸��d��r�n�^s�����=*�XF���iܕ�=�-��_e~G��Wb�ܧ��֫��8�>���6���!��x��=��#�
񯯘g���e򞏜���$z�}�w��n��ջ}�˩�U�*N�rP�\���M���:��JXOݗ=W���2�a�Ae�l��Ǯ��pft�Y%R~-�=Xq%�����w�y�KnX�F`����cp{&�>�o6�joܶ���Ӌh�,�ܔ�Q��i�S^m�WI���N@V��'�?RG9|�_�����x��x�n[���py������`ƈ��h$��j��z�p<Xy�B[[��h�=yW����X�$�F��)G�hp����aEvp��ہ�o��'6"�!���rӷ�*}u�ѻ�Xߦ/bt��K��pd�@�mڢς�am6lL^���௒�V"��̽@��d�Ћ��T9�Yñg��ќ�a?���k|l��#1a	�t!��J�:�40�sV5%���y�X�)j�<��TQg�♢�x��#��]�(^>!//u=�b���a)�S1��97T�|�<���=�<��!��9 �z>��e���x~�Tp�<*h��_��������2��T�*z���h=����J\���Ip�� !&��Bu�5#�x�3�aO�'.�|x�ݗ���������zhX�Y���ѿ�@���x�Qc^)��R���yN6�*�<�t������(_Y�5Ԓo�y>4���羸���������I9�_H;��WJ9�(�_tS������Z��4F����)��z��g���n����/n�fۇr�n�	i>$>��2�\� �����w�����ó�gUT?崷������kTGu�|<`�(��6�0(gr��/�E<;���
���ZbCZ��56�竢��CE)�Q+̟�i�aM�+�ƈpp1��I���(�	�h,L�ؐ�(MbU�0�v�4�ޭ��Z^���6������i�R.n��p(�*&fwJhs�$V7�p����ц���6YN��y�:9��w~�p�Y��2�i���Ɇ"��+�ߩ�]/�Q�VYY����[�'�~��xFB4��W��˩h�E�W��R5)��rY+�4H�1ՠ	�i��k$��Y?�%y�|l���h����݇2�j�\�F��+v���;��r��%�1�6��N9G~1�C1d;�k��A�O#����a6���e�����}Y�2�<8� ��#�c��8l2����x b����D6��Q@��� 2���N(jh�}���=Ћ��۸7�X�s�=x�x��t�'�&/��S�Mw�cP�|��g�
���Ǐ>ִ_^����'�{�Û�x��axp�
+Hgc.C�1���ށ�0%I��n߂������g1(���Fј����^&:�˹�f	o��GA��G�m�«��&|V�`�b��N?���|�ku�~��FŅ���,V����j,�#�GZ1v�ሊ��?3�^���^�*Wn1?��V�d%��4 y�b.Gc�q�
8�8W��R�l�~�K�ʼѷ����]�%����AO_��T��с^���B$*4��7�����5(FF�׈шa��?~��p9=�����"��h]��|r8�b ��	��������l���2��S9��_)h��FzG�g��HJI��u4 4��t��)�
�oh��P�=t�E��?Ea��N�D��>�=����lz= 	$�������̥ؾu�za��0�ƪ*(��Tz�q=rKm����!�Q�P�Ĕ����T4���T�0�i�(�
ܴ����G�gO
��)�j��k��CS2=��/}�"%�\S#�x��B�utD�*�Y�MD/�J���
��2eUcC�&�<���Ba����x��s�1���
��Jj��c�у�҂�p�ʗ�Fݜ��(����n��](�\��]��3v����lW��|݋����	YrV�e�����%�ݺ��N.$�����Kr���J6VPAɡ7�um����M����z��k�L�{��4
�Q��b�w����f����q=�]*g����i�=Gs!���g"�eDb5�J_�i$�d�x��z��jk����8��@�m(c��C�:�4ܗ������HFC��Bu"e��1rq�q�Xl%�U��"9���6�b�ce$("����=���Pgs@���z8�q�SY%��&�Z�pod;���,��� ��(���e������dVJ�'�rj[�Ѷƃ�Ƀ��T�V���@x/tm���VJ�<�A�vJUg��[�Y����ߡmmc���\������y(�o@Ձ�w��	�o�4KjԷ���!`���%Z�j��lS$�W6�Rӻ�1��3h4���Y��&����O��8vw��x<�Tx���~�L��f��XK���Q�Z�Ե��J7.�7]���w�,G���st���Eh�U>�SY~���W�`=�HL�w؊�[���t���(a'!�ˑ��aK;���Qј�Լ]�:��:8<�P�b��e���Q���X�X��e���2�P�����g!*�8x�P"���E2h+V[i���e3������<�P�
�����o~�u���<I͵��T�^��\��V2y�ǜ������+C=j��A4Gq���^�˩�����o�$T���/�Q,�&�����F�.qs��ۈIncy�FB~���]�a-�����ШH�j�.�a��ǫ��
vʰw ��:8T�*V�Հ��ew���6�ω8�iY�औ�ށ�2��y����R���<4����z@�2mfG�p �W��~����ߦ_��^yK��M��ʡ��k�ʨ�(H���CQ�p�L�n�*��o��$a�"�n�d������=�2��a�\������Ո��3����<v��-��f��۠o�B�o5A�@nc�|B���#��8F�W���Ÿ��=h�W �;G4Q����R�v��j1\=s6|s�V��G��ճ^_�҇��@G/�U�
oĈ%��:1�� *�����a�ư�1h�Q���L���n�Q�*��m��{3Z�Bsw�����E*ĵB�%v����Û�P1	
X�A���&�3Bu��G9~���nXw;)�5�0��c����jT�N�ˡ��o��}����f�7�X��|�!b�D6�ՓC.Y������7		�HT��P�X�y�9�<��F=|���T�:*w�Q�͞&�52n�߅�������8��ĺ��K��q�����mk(���&�U�і�|[�R6b1�Q�F;.���2^�} �oe�|�������0�-��r�CʯwVu��uҥQ�˵p��q�������d�L~��p�qf�,�o�m�x@�t���g==A�+@ıЀ6Z���o	$ÁW�;�&�ǹ���0�r��������6obrY=%l ��j<i9�0$}�#-�/��+�T�9li':�����C=��ֱ�r�ny��h�m��<��ԉR,��ك����^�+ڈ<�y0%?<t�`T�[���?ʼHmn-��̑4,�w���W~�`&����m�.����&9��L�pH�}H>�v��>X');�x�*�A��֠ )0v7�'waE��wt�P�^؎����B��X[w��E�/�qF�<V����s{o�R���s����=��Tb�����Lb
��t	Ǳ�ʪzr��<Լt����$�N��N��؎����9����ٱe	��B+�m���^p|���gn޼��
WH�Ν��;7�H���-9���5,	a%��1���WfVQ�z�x�D".��WF'� ��m��J��h�<N������^�Ic`����=�c�a��oBP9-��Hiyi=	��Vp-.^��2���a�`B��ÎY/�N���t�_7�݄̳*;���y6&'�*��{�ŧŕ8B�ޙ�}�{Q�̞�iҨ�J�I}d��h8j�[c�D	$Á��
���%�y?L��ƍ^�� 	֍(�en��jA�X���Q-� �kZZ_]��R�M>�yuu���#�o�dSs��Yl����G�����������\,n6���]�C�Jg����f�RI�Nc!R~4�%�7�9`
�Ip#���5yL�M�N��=B.��Sѻ]���F��\�z3b��l �i�P�OރP�<dsx(���K]������&ɝ���KdB^����(�ň 皺Wɯ�b�v<���b-&[���=��M1n^yN�)�ѫ��j#���'g��=&q��������ब?����Qޏ�3�>�2�>2b:	�E��/<�S�Y��q����=�k>��d��A%&D�Jo��2i}�b!-��˨�U�y^BC 5��/�������F�'���;a#��a�Z(��9���^z)�J)#��z�<�I%�3���=κ`#��1	sI|iN�$��\�`�A�z��G����Ͼ<�����P���*d��y��$����(�o����~�*�x܌V����k-p��\/s7�{���3��p<(���<��'Ȣ�W6VV_�l�s�xT<8�j2�n�%��y�7��qc�k<�M�����~o�ʁ�'*�CXF���[(�L����x����͍��Rmes�\�h����4��K�19�zQH����5w2��(����S���y�P��hދ���fi�@����d ��R%,߾���~Xa(S	E�8�\j=m7(Ņ�iz݌���[{�5Ob�u`$�b螑�ж��.��>�X8s�L��]#��ΝB)����UF�(م6�Sv��6Ʃ�	�*�<*� G��JV>����P�W�)�$�rD�2�Xe�l�aT`F����b�����jF~X1���we2�u���`X�z0�F�ek����Zvx3˙1�I��6PnA<�63БpfD<.��x	%<��-���JVYaD�9�M�TjoOOw�A��Uc�Bm2+^�gz2�XWq�('�k��8#PV��+4��N��;��o��hP�G���3B�W�۟��x�G���F��������@����>�T��d��*�$�-�1Zp]�E�W�9�wn��d�̦��^����k��젠bc9|�OQ�|��m<����DD�֖�,Q_,f������RƘ{·��W��XG�Wk�!��p�J��ޅӲ�J�~��n!��Md2����
����o!���[aP��C�خ��cS[�Z�46��wJ�����x;�p�s�)'՝�1�g��5� ז�nR���f�����V�y�Y}�W;3���������f��x��ez��-&�x+�Еxlm�p��'��/~/̭���g?�w.<�p�1����VQ�Lt�ć�{�EZ���S����ݳ+L��ƀ�7�����P4]D;z�z�c�gVHdG/e����W��^�WH5�82��8(H���2
����qE�e�x(^�ܗ����7�S��by�N������[+;�rT��Te�������<����Dh*K����{��$�j�l3w!���cF:%�J�`���.ܧJ�~=~��1�x>�'�mt�_�3����m��m�3��0X�k�¼���ф�k��A01�/�TN���p���^h,�ʙ����mh�ܷ��y�F<L�J��m�=�5����h(�G)�+4�~{o���]3�y�@�#�؂����9¬��y+����2+cD;�^#�)ao_��x���g7�����7y��p|�n����R��d~�7=>h|���������� ��e����;l�����x��0σ��4:|�p�M\[$��Jv<�:ɛ��6`0�ٻa��dx�S��������x�[��o^���}WQN�$%��짡>Y��tu�ļF���ڨóE!R�5�c <��btQ�Q���TBBW95��ê�Lyg�U���
�0$֎w��QA�g9�����r6G��iH�n�;͆K�]�*�ə�u*����r�,�b�>��f���4q~fᑬ������s���Uw�$y����R��7��6��4W#�y��s������Xr*D���Yo���4��eܿy?KWbR�++�{/����~R!+e붌R�H4r9��y�O9��M����x�CxL���ga���p��
�jf8��EM��� �;��"���5���Xj~h6�l��{���a�Ȥ�@�%��5Jo��2m�������,��n{�%���R����l���T�����gŜ��Ǭ�X��(���}5��zxP�w"�i<� �Sי�w�z8s&\�@��ֹ���y5\�^	�]aH�['Ù����������_�Je(b�+�A�<��TZْh��Dp��MTUHҏ0R���;*������=K����@yZ���*+���M��Y.��"L#�G0iM$bC���-����˒���j�C���yU����<m��ȱ9v�GV���1ۂ=8�R��s��{�_$e̍������y�2��ѕrX$�R����U`Ng̍��D�Q&RYkt�<v��	g���vdI�o���x�y>�#�U����q9���?ܟo�w�V9���CH��կ�(�}iH�?��aR	[Q���x�8<�8ۛ��{��^��sF]y���;�F9;΁Fž��`�F��ؙ��yͦ(��̢�"2�eܙp U�UO��4�O�Zy��b�X*6*-�6���@2H�����ֶUF��6
O�36ϡL|P5&���5G���ب�Z�<}ԓ�φg?��Ѐ�c�aPS��~����]�������������e�L�!i��yhg���t�Fx�ӟ�]�R�H��j��:ǂ���]'�br�"�)�&�����r_��i0�h��)�'�9cEm�V�:/����BAQeH��?\7���ąy]+L�OZX�F8��ZVa�j���e.���ʌS��nD���J���@D�d�e����P����6�m�x����-aՀZj�T>��߽~�/�,��rp���rfR��E����_��|�k_��%���s�3��ȅ���
���hu1h�,�5"�{���v�oM��e����M#b�%���x=.)�5Z��߽o=��5Em����xy��Y>)�6�\���UZ�ʥf*ȎƊ2!],�t��Ӏ��Q�3��OLLvsLc��uV�p|�������0�5��&f�)�U *_Ǹ:�N"w���%l���p�Ï?�@I<���pT�D/�ø���̐�`{�7ަ�p�~��.�Խ���/�y(�wd�����C�*�.���7����㩒����é�Ø߈��$��m�1Lc$��W�d|�9"�L��G��`&��0�d��1�?�'�y��B����ik��kR2�˨��
Nn^m����2�<w�A��lNĭd0��cՖ/=����ؕmC���:�"���L��xU�~��U���&���BFz��j����پ�F�y ��^�Pã�5Q���(�o��/9�����/�s�������2�bb�V/=F)�T--���=���^��{5�%��pl;q�)�0�����������׹�C��+�q?,���<�"���K#��4�29�����Ժ��ҽ�p�Lz=	$A>)��6����ѽ�%3E���l^�tT&>�V����x\��*�n"�u������݇�� �G)/F ��Dޢ�~�%�u�7�l"_r���l�������9��.�	g�3֖����������
F�Z� T��S��}$�#b�[�&��V'�hχT���r̨��8c��qNe���I�"_31)�S�Њ�;yS�
9R~�a����5J�l�4/�4�����!)��("��?,͠�X����s�ǹ�Gx��}��'�W	OO�FřQwLG������#��1��6��ZQ�y?�����|UF���^�g����4Xn�w�G��0
�(��]&�qx�܆���Ů���FE�g$�:�?�.4bBnVbY�m��$7��^1+T��Lƹs�*7���J:�v��Ή�u���������F3��>���#�� 9�Ǐq��q���r����$�"YH�і�ɥ׃�@2B������� ���C�7�	3�`0Tb�> ~��矞��压�$L3i��`����Xo�t��$n�I"q���$�5fZ�?�b����?A��U�i�B#c+�Y�p4��81I	j-z�x��������¥F1���9ŉ~$�stT>�[P"&�Q�۵�$(4&�U���a��4�����{�~_�~h���mdQ��Ի4
���a�hq���@t&Q��C__BL��Y
�G��"�������Go�ٿc5�i٪�^��"��ڎ�F~��w9#�i>�Ug o�3�P�BO.���Rϛ�������归��u����6��/��mh�40�K���C9�x�����l7��O���"��yj�5�{vS�l���<Z?�h�F#���̳��D�U�V�Ƣ3�]���OC8�B}�"e�L���FC��"9�}��¬�.#?;9�&�+�@�����SW�'��y?�!���CީḂ
�d����,��� uJo�<�r�����53���uF��I��Ed2	���?�>�N4�k�� [�-�jh/��7�Cax⭒)���^�3=s�lLBwc����0Xe����l
}�D�
Ee��jTRn�����;�j*)�vND���r*Y�[��Ä�	Zv�`�U�U��J���� � � ��Dy�)A���<�ڪ�5< �\�[�J�\�� E�)���QO��Uj*Ϝ�=K��ӑ}���f^����ܶ
��f�-�������e����йN>
V�\�(!��bv��"]��W�F���
Y��rw?��2b�X��� =��F�ur�ssٜ]�c��s��hä���w3Ӕ��*�\_�k(5ZB��*7��܀���Y����l����N��YV�]�5�C|��NDcQh��wI�L�;�w���t4�i����8�~�Ӵ�GH��cp7�@m�$�
1�pۇ�h�8 /@п#[����Fe2D��n��+z��8���
GQ=x( M�Co1q�r�.��8��Z��2����Z h� �iw@�L�c�v��mJ�S�9G���=*�5��-`�i�җf_{�V��M>���L�G�A"�H���<��4����I�We����9���
��T�Bp������Sx����k> u|sG,Ǽs�VT8BT&ȭfc�z�\�1�.ǲ��C��|�ƾ��:�H"o�'�"���g+Ŀ�p�:�mZ��q���CE�{�*r#
=q�<G�S�kh�:܆�o٬Jވ�(���گ�Z<v#��	�M�۾)8�*�O>�D�a�� �%��3]�-�AC��2�)p{V~�����2�G5H�hF���zͯQh�_���[fxk�1���q�>��w�Y%٥�����4?�p4$'���5��Q�:���{�s���T�̸�ʱ�����>|��䇐�����8E�ۖ��K^c�B�Y[�x�L
��B3�I�ϑ7�p��fo�2���xt�mЛ7m���a�S���h����>��P`�ՕE���PX������I �_��߈�W���
r���m�H�T���T��p]V��wQqD�ӬCڷ�.�T63�y�����*<��+^���co}!���>�
2Ш|��XƑ�sQ���KڈV�]����ѡY3��z����!���]In@3���9�aeՇI��y��2���5h*K�b'&2��|t���R*Y������(EŬ�T� t����_�|�
��e4�2��.$��Lihܷ��x���o��{.��r1�Q2B���u<�<r��;6�4b�8i 5*n�*s�G�n�{�m�u��Y�����a�{��FJ�&���n�A��hԩ,E�ҳ7�(�)�W�8�u���J<�h�LD�����/������C�cs"�b�����R����}l���k��ܼ� J�_><*����||6Q�2����q���0�\�><�8u��6�����dx��������]���4/<����p�J�"0�[�槫q�:<T�������q��3̗������������(e�f��:3�Pĭ)�WPh(�A&�|�f�a���ؕL~��W�SɔsW�w �*�S/2�DF"$"�cY�0�d'���(�
���9�� �?8��yu�o�<��޵'��iGX+Ν �2gD�UKG��pK��|M�jL��1���z#oV�N2V�,q����Df-l��2Q�Z���ԓ��F�9[��飊ZÐ'��~��mMB��P�jl5���k/,�×&�-��8j ��m,����A�eD߸.�6�)1Z��Hh�̻x\F�����j�ܶÿ9��7z�����P\L�_��[4��C�=&�wzb2�q��L^-F�@M1U�͕�+�4t���9��
��&C	qK҅�q��4J���Z����tF2k�� ��K\��3�o��)���x��`�Qh�G)k��ҋ���[���6�lt�k��;,��_�hA�u�>�����V�ͯ}%�ql�� �� �a�	�!��x�t�8�������Nc��������G�}��9}�\���R�w2�iü	�P��3��:]�w��|8-N�3�A��Z�e9��!���"�q2�ʢ���Z�	���[�_����G�x�����cy�^�72�V�����
���nj�r9�^�����ǲѝ[��{u���� �K�AV'p,Fy����{���F���ގ�x��0
�?B�E���rX#�%����8�o��@e�v%D4���I�Ze�o|#FBKyՔ��d�/��{�4�@��$NԸĆ:�Г�B�dt"D�o"�z�����y�(��7C�%��e ����ԗ���!U�m�"�mp�CF%�}�F��\{�G��79.̥L�����n��i�}r���J�%�q�#ɭ��ʠ���ޛ[v_�}�;�;Ϸ�	��n��A@�(QiJ�K���q�$U.+Q��T��g��خ8e���eI�dq�Hq Ep A�1=���}�y���ٍ%��@����PWݸ}�>�|g�5~�[]]ˆ����^ɛ��hi�BCo����֘Ih4X�Ǫ>�`nHTt7�fڹ��P �������::V�a�6�`��F����!ol��`� 7Z���J�}4�)�xC�2oR�d�0�����mAjb�ʵQ�_'���+��;���!r׮�dc���?WP$����X���H�O�)sg�D�2����3��˂(> ��f?�憡:B���O�Lف��
['ɥo�W[	Iv�Y�i5Or�J>�������o3g�]>ETr�A��A��ce���3��%%�~��a�[������a0?�3+����[d�a`wmۍQ�A�v,��<|o����iX���^v��05� ݞ?[���r�����q;���y���ߍX\U;&�%������D6Eg�y�y��,�>VM�ՁԚOuYI�±k7�-���P� <��m/Ň�R��c�O�P-�n��­�#yI=��g�{>^�:����H��^�V|���Jg���'D�i̐�,���i��B��:�%�5��\��(�賝8{M��r�١�0��<%n�0�_ 9�Ğ�m�s'����������;�*�I�P���q�)8����#\��O��A��	V�qn�Yn�����co������ů�-:m��ӓ���r��8r?���Fځ�؏���Kԡg�y&�k�w��竔��h�-l,��: ����6��f{�E-��ɨ=���N�m����oŐ�3��"\���<�ͦ��o�@V2��&�c}(S��H��ϭ�Da�_�3l�3#�������#���r��ɭ�⒢;�y�<w�Rt�a��a�1����G~%��o�Ghd^���9u9L�q]Z�&��i����uP�͡�0�v��X&��B�k�WK�j�(?�����|��]G�h2"���cWo1�b��XTx�*3��I$M�Q��f]��K0��v�.��B�{���zI:T���+���KM2�����`q��\Pse0V���`����s����}/_�s�U���}�k_��QMg=,5y�u���:��AX���kG����j������{{�����1�oS��k�T=�v_���Y'D��	�*�5ٝ��
����<23cds�=~oy��iV��6PN�����{�[y�ˇ�z��ݸjś���溺���Jַ��A��z������峃�<�̯3���m�>n�%"�yn���	Ewk�o�,��elp37��;��Q�(!8�����7��f����6��R�,7Y�i��3����y���!n�ү��b`��7s=�\7T��������7�W����S*D�(�,������7�1~�*K�'�C\.?��O��w�}4�����ë��
�g��0Fe�-�Q_���L���b��4q���̶l�	34ԕHim팈YCV7�urFÖ\�a8�o$�j�d� �%-����W��A��)u1�?��_5���=0�:�Y�q��CO~ >��?���/��oF�X��Z���g"*�`w9��J��X9�'�6��03x�!���.�Uf��?�}�؍ȗi���*��aȤVpʊjx-!�f�#�g�}62ːN���9eH�,,?�Y��G֙�"���I��ļ�D�H�$tR:�Wf$b(>�_xl�nVciM��=��cֻ9�m�.����{����s�����������Tg��	Ճ�������K�2�8��nq������-��¥+e7=��T�6��{�~�~���75�*���Y�mǶ2΄yw?�&m��܊~B����?�=���VF��zP���k��طu��Ǟz���y��G�{}unepses�m�m�?��'f�g�W����������e�Ƙ��ʟ����P؆Ci�}��=�D����o6Ʈ^���Y_eGY��k������sv�m�������z�N$}�,a���7��oP˟�O����.���ZL���Qz����;�|�ll?\N��,�nRX���Q��2���&�;ï�)zs���å�PYa?Fǀj���`n�xޤDԹB�z�
�*�ew&@y,�l�9?�t�Ϸ�F�|�&�-,}�|��
�Ul�[v2���2���{���]�r��C���5�#���{����-��X��Fõ97��E�zv�W��~Y�@4�����>6Nݜf r�L���{�����Ksߞ˺�*��-���'�N����͆<�ŔFԮr@W 0����>(r��s�0�Ȇ���Q|����#[k�q�]4�m�+wϒl�m����{�Ⱥ+�^QN�i��#��e��念����Ev5�>�Ç����ؾck0�����ivs�w����)���$����[G���K��s13�ܤr�{C�3(w�r�Qs��q10�W�q�zZ\_-���1�d��'>��r�'�m=eq�l�?����fd��7�"����W�/[�aU�&)��f�S@e�kg�����(���R���ًE�����v��Ο.�lx��z�+o+�#���*v�l����rٲmg��H��?��B�5��͗��(q�s���T�N[џ����gC��;���{���=�C��2�e�1�������$~��h���ǣee�Ŕkk��`�l�u}�^���T��A"�D�kD�X��q��Dj{�.(W|��������RO������s_3MD�ʋL�N�㛾C�v��e���y����?v�`�v��5�菽�J�V�F����81;�4�@��v�:^�w�R*�,o�8��G���g�A�y��l���,���1Te�G�"JI��؍p�W]�4��˙�ll銨��<��(M��),��0��MV�Wkv�:�頄��n��ęlۆ[`�����wk1T��s��g?�����G>��1oWy���ʃ�WF���kWΖ�4��o�IY�|D��b6ס�����wOWs Q����R���t<�H��3��?���$վ�&E7Bћ3K9���=���IJfb|i33�JfE2�jE[���mK�o�/~f
F�ʌ�=XZ2K1��W��D�y���c�*��@�����,������/hؼ�Ƿ$�j�.����	��i�1�s��Ub���	ќx��>�ԙ�5۲�e?�&+�� ��y�am��P^�ɵ Ӭg����{�-��)�dW��?�d�޷���=�����/#=rO����v��IH6����7U�9���;�����������_��+�_��h�����u�vi��K�������������k:m�#1�a����1�_fg�[�;[m^/R��=��6�-�S��f��ǉ,C�\cN�-}�G1 h"�����������=�G�.h�_?�(|�2�v:/�"�VJ
�����u��`�:�ue�%2�j0+n�`�V�{U)���������_ *߂��;N	c��
����42��W�:(H`#�G��a�C]{�5�D�:G�G������uF:���b?�ё�s?�hd����ֳ߅��&�ko�ZdC�9�ʥ���-�Sr�#�a|�=��4	iu>���u����}�J?�.g�B|���ט(]"��zT�	�E���yA��8s�����`s��ɷ?�S��Dtu�[� v��|�Y�s"6�=�eL��"�0�,��}���z������U����秚��yT�E�a�b#^P�8CK����0��&]Y����M�Qr�:�>�ב*��7�'[a�@ז&�o���J=�ko��z�Iط�ٻ�*��sK��E��4��tД?w�by�`���&ExQ���p�:�������� �8�${G�)�w�ز}�+ioX�s��;߲��,u�K`1WQMs=���]b��.2���X��q����O$?��:������{H���i�J9�С����=�D���A㱋>�$5�sԏO_�Yf�a��XBr�NFK��Abom!<���O��5�,���t#_휂=��4L�1�jZ$�����`�9��8pC4�ݥ��2%�m��>��������Zl.O�X6q����i�X-������2CuG°��3T>����^�Z�<���]��S��L���w(��:�v��g���T5x��̨�
�Ѿ5�G/��*�:�מ�5|M^^+[L��SδŘ�y�������/=��^{�͐(qˠߏ���%�B������k�H{��I����YU*�J�}�7cū_�)�����w�D��͌����쩳����iH�0��XVCe��ƚ����g/�f�q�&EW�R
�`�9�aR�1gE���kG�Y;�a��}^��qy&���rݴ�EzI\f�:Tzߐ.�Cr��镡�FV���|�r�P��]�R6�oG"�ѲV�&7ÿwp/�K�,?�=���A}{~iqu�]ئ��C�K��*�[�F"9�{���0K��}��HZ�@�Է2��J�^z�o}�_����`�C��A�w�{غ�=s�|������2Ǎ��V�"��:NC�4������5^��ȝ���ڽk{H��/�V�D�����}�J)F��d�,�vCw�$��?9�0�d�͂���P�PXQ%['��8vP{����Y�Ât�W���gm(tM�C>����L��/M򚍐��<�	#�ԙ�1n'��;���X�Mv�Lc]�j踣<G�^�����j)itM�O�������P�%?���~�\RT5�nųo�t����Q\5��I��I�cpV��_���e�]���c�:��6z ׯC�%#�A+yb�P��λ��y~oY̞���5a�cS�A�=D�/�x$��:�G}|v#�zc��ʌG'�g��,_��I�*[ɘ��g��^)ݺ�K�B[���#�C!�>���Q���(�P�z?Ô;ɼw�t��P8!?�ߍ�����:�ƉXz�E�`��^�λض�eC��B`�t�����d�q'P|��`��Y���.��K���ü���ODT9���$ϐ�؀Y��B�D�F_�-��ǟ,�O ��8]��@��/���z%�Ǎv���g.]+�=]nP
Xo�����E;�8�+Qb�os%��Y���cǰ��tēO<^�y�5��N%ҿ����Ӭ�q�%��X��G�Gc�ǌ�"�ߡ�r/��z߃�O'�Kyng��>fS:i /S���PuZ�o�X�p���Kd?$¾�^Go��O~����)V����ۆ��H�H]@�� ��=�1��hu�̭!�24�i8�P�U-_e;�m+P���wT��B �6�俯��iH6�=~H}�-�L�=1>S���J��3g��Pv�����|c�of���?<rf&:�m�J:�����n�D{ �2t4���{�	��c�IMs�c��C�3�����<�8Dԛg)%z��b��e����IiM��DU�:͸6qv��eM���v��:�:02Zf`�y�Xۃ4�3��X�+�o'�#rI���>Ts}��ɪ�AZ}�2<:��At�d��6����Xj����;�@fw�ww�����S��5�!��L�̨xێ]�`�Y�pj4�b�x��Ѹ��s�J�/Q~���w?�X��'�L�\����^���O��������_�z��+�ʕit�`�4�o�C���(m�����:��R���,���t�A���$��Z���;��r��j��;����6C�b�i�b5,Q�{�[�s���Mh��4�y�}D�]1��<���Ns|q�O��KU�z��t���e0���Ç�.裏����8@Gh���ū�jŨ����`�-���E�eVCa,S�V��*���Ϡ�_g��U4�����3rW���AI�딬���W=��ٯ�<PkP�%H��dO��W��u
5Sʷ��/���n�t~��N����K�4����s�=��A�]���ˈ>�+QA�`�1T\����y��
N���XIw���l���ۨ��n�ņCԉ4�3�񝵀�*��3_�L0�3��:{y�k	�{dܯ"�A�o��D�����7_����DhV*mG>D�$�{l�����"�ww��+�q���Vv`6�Z�d<ycȪbz�r�7���PX��_�h�oi��d�,�~g��F�ԗ���.{�{�|��W��YJ:C{�dQ|3m}��I�F7]?mDn�e��(�X~�&�5L��wv�q�6���ր�fXt�YC��,�RJ��/��Ғ�L"�mFӖ���W�>y4�W�����Ә��F�h��wR�v]��а66�u���o���S'ϕ/}�p ������(YXAn�<j��nXkH�\@�oΒ���\t��L�c�7V�6��q�4{o3��RU����x2��f����[F�6�癏��:�n�..�d}=`3C$���,�x�5d��\����j��N�8���&e�/|�վ
�Ω^��p����:G�	��׽�Q���tT:3�~��+�W���S�;Ġv:"_/�!����t�u�.03[YQZjj}��X
t�od;4jcd�Sseja��s��K�0�	��{�g@?�/��Av�;|����G�B�R/�0��5SAP�� �1����xǽ����xϝB:���WB�vuan�M�/t�Im�q�%�Ћ����@ҁ��8�
�`�̎_��L����b{����k����/�;��m,=��Z�{F��TC;��,z5`��~��#�}�p����A��V�
7�=R=�'�I#j4UJ;!k�+��48��[0��,54���k�ltz��D��ѵ�f��f�>G�~?&�-�`4��$�QM�6�zF�:������~��c��)$*6���a�X��m4��ʹ(�){b��*Q���s0�!��t�"�h��Y_��R����F��E��S{�N�Q�i��!��z7�6zPw���2�N���=�Ed\�{�;d��yx�fJQ��b6�����+f=�3!�q�}H��y���g�^�?�|��8.��=t�������{T�U�ލ����D�p�Mua3h�i����l�:�ܫ�o�ȶ��>_���mr��ٌ6�O��%�s;q�o��r�a�ѣ��˜Bߧ�?}
F;d�<�b%���N�|H�^ь�����?�SH���7���-�#TQB9�)L�a�o�������c���|�H/a_V"��N��@V��}�uxw��yw�}w��QZ�ir&����5�A}7p jXiH��{�w�r
���rn>"q���q���7��oM$�<�~�i-]��W��eG��5��))��~����=U�i�wb�?+ʕ���kx}el�Cv�s�j��jA�� }�ӭ�|�yJx����O¥G��&�T���iq��	�G_og0��b�z?�l#57J(��S����[�hk,+�?�̾�D:3��s����R����6����h�<�M24�t~�(�EP!�F�Y��z���y�ODII��13��ޕ;֝"WWʞ��r��A��� =/W}{~{Q 8t�p4�u !u��@�LH��{M7��9��W���ǁ�=��f�:�%�Rh#s��9�+PM�V��.����K�3:TE��c�E�*1@��Cn\<W8�`$M�n�s�!���|�+d��8�[�a�!��o��JV��H��JVW��������B�W�#*���*��1�L�a�l�ފ�Ĭ���n��[��l^-{�(W`��}�=�7�$��Ϸ���GD�A��.��C�ԇ�I:j7i��f�0��D��ބ�!�W�sd�=���v�D�d�v���T�+OQ��a�K���t�LȨyz���o����aO]��w�?��B2���Y%t��3��[��ဠ�ڭ��N��!���-=��8�=,���y����~�|���*/\-�����,�kt�ܜ�Ft�;jg�"��������.F�y������L�?����
j��Jq[���K8q�eD��C����f ͽ<;�(�h%��[�G%U�q�ﮢ�VR�f�β�}��m�[��a��G��*#[�k߁虘A<��Q�b�I]����]��ػ��90'�tx�v�X��dI՟3������7w��;�+Z��T�Zb�U�Z�#�P�	X���B�Y��GO��N�&U4Z�v"S���>@00S��}��/�Hp��p���A����� S'�������o�^�x��쥩kfF�t�*Og�����_��tw�wz($��0�yUr|S����;�:����?K]���sS�_8Q��&/O�Xb�ƴ�\E�*���Fh��|�E�q�lQP$�n�8b��"70d�%�F7��t�h���V���Yf�`�9�GV����iūy�1�aI��\[�(�Eo��{�7��3�;�ul�'24�1b�/��lȆ��Mv͛u��WwL;\�Q�Lч��$e�嵖r�UÇ�w�%������o��oE��o�I��_�u���p;{q�F��ϧ�z�����3}�*�A�zh��G󀇻;����tSNF���V�L(�wҌ�i�ɀ_���1��Neu�H3���݈:�=��x��yޖ�T荽#d�]Ȏ�����x̠�^���5Qɠ�E�3Ky*�Y��I�e�+�O1E_����W�	)E�@L>xnt���p�Я��z	*�1��0�Ȳ��<+`O���kx�~�52����ZP��L���X9�}g1�:�� tA�>���$N�K��;e��~��׫d�;��:N��& ɱ��������y���
VPqd�D?�� o\n�)7�q�mN�(�y��^�P�./�k�e�&ƏH|}�}Y;y�lL��Yd66gip���}��ee�:��,��}���E'����73Q�u�%��2^4�NF�`8-��y�@���Z5�s!��,�7j�d�)n�az���Q4J���D��!�:	̿���R���snR�۱�.j�,0B��?��7Jr1�'��ـv�|���*���ύ]��w7�m����/���O�/��8T��~���ݣd4�_}�7ü�R;z�L4������Բ&�mtX�d�5�L��T���ԫ��۔S���t|��p�#�lU:�%�x;��㉗F�L@&���3^6��.�Qn3�����`�kt�U�dt�ϕ%5���j�}�s)���j�X���g��ݸ�|1ˊOpk���K�T,MVΦ��P?+
߅?k:1���:�����`�u(�9����/1��1�\�����ԥ�em�j�E��3��_���m���������ȎtQ�t�b8��5�X��:��qm]fw�wz�����/f�Ee|��z�!a��1Ճʊ������߃q)���n"B�T�F���ͬ�*��6n�$i}�A|*��u����X^�����ZG��PX�r�b#�0�7�=�r�:W��[�n/�2�.�Dt>O9J��K��y�Y�
�2�M��\6C�~�!��O`��Ȥ�l��)L�O�-�u�A�C��_���D�a��X�d9F��>�w���k�>����$v�#O\~��Xv��uh��U9���O����2�r���/"Q�\(��k��Y�VzlE���F�ܣ5�wNh��^DDזo�;<bG)�ӿ�B��,w
��ԫ�Fҳ�X����5辧�b�ߩ{!:�(J?�ɛ��x�A���ۛ�:wQ��<_3�#�/l����a*�1{YM'R;�܋�>K]ʪg[t����~�e�k*HZl��p �dB����j�;u��H�f��0-Mm��z�.�Ɏ�ۿ��{�2:�R'�gwɻ�f�`�4d�%2�1w�PRl�Ȼ��ʊ��-�©��*YÕ۠A��;5P���q�A0���q��-[���qxI	�Ut�z���˃���!�Mt>�d-��>7����3�<g.��������uޘF�m�Uh��8%�TC��amc���C}�72��:D#H��j����5���>�N����N*��Ӹ%706`����9N��P���d��,�B0��'�b�D�l�,Hè዁<����2��ët ΦtE�s�Rg9
4ұ��u��L!_�����_�����i039��r����O](/�Й�\���7f#4�@���8�@e��j9H�g�||,���Q�s\0�[��0��_-�T} �H�&�8V����0�M���}{S]c�Q�-�����Nb^�y>_����2+fΉ�{�!�B%�b�����y딂� 3��ح��vQoG���/S��S�0�K�`���,� (�4x��J��ܽr������ C,�!H7��� �����<����?��(Iu�,9�\�!�^�,�=I�y�����O�<kLq8W]�$���_�[����C ����;?(�c�5.1XK��r�02#?����O|�Qd�i����2J�i��p�9��[���E�p���O'��Z9~�R�y�|��}���(��~&�or��t4��k�O����~˺�w�¼���GU�F�W��c�x��*:�?q%^W۶����G_���{\��]��)�SFY���4I�:�����_���F�fC�C�N5'֫&-烌��8������������[�l+��݇�I��'�;���P~}����Q��>��FC�c�R�����'�@KU�C�dD_;�FJ1��[c��c�K\����&�*J��\jٖ`���hR{;�!W�%3 w���Wa�5��2���0���,3��)�>���V�VY������^bUS��rf�,�bm̨H%��v�r��|F��j���@d�<���'Jf�&C�9����*�q�2��8��ej}�\���>���_�;�k� 
���V�颼������� ;P�!Q���^�a>X>��)GO�Z?WڇF�_5Cƫf՗���㝛�?��tw�wz��-=s=k-�Ԁ��v�ߡ�};�Z����S�cއ�[�M0���Z�爦֨)O��1����F~���N�7^~������兗����`Z��Qh�S[�.�D��g\��]v�^��7��.��֢��V��C9�;O='��~��6N ���x/D�:��'A/�lC��4�H��:K��f�h��ڴ�O��)>S%�.z1���t嫯�!���A�p� ����:4�kD���p KD�(��M'��~�ָ���/�3�}����*]k�U�:�LY��F933=�q����v����J^��ʥI��K�{C�x��0�Ȧ�γ�gn�`��=M�.(����O�88��V��#�}(
7�W���P�uunlW�8���m��gm����|�m�t��tP���3o�K$6h�1�vk� VD߂r��18��`��!;O&�����Ɯ�*�fW>��h%#�=���2�׉�7pAWKe���k�iR����K3k���:�"
�� B�rqs�9��҂��g?���S��rh߀'-��}2�x�5)zX�mVܿ�2�_�d��7�<�|�nʒ�Ej��������9�֖���2R���qGH�qG`|w!B\�g}�����0�7��~�s���^��%�U��������i���ж��!}7�˭I��Ð7�^x���-/�q�����M�w�v��Z�T$u�S�;
s:C��^�u��*#��[w�� -a�1p8Em�.p�[�*\uv��P�izz>�u(�nʉ�Y��A2�Z��.��a��U�U��*���Σ6���9+PQ���Rbt� X2r(�[�� ��'}������ؿ��g�zF�ly���c��#�6�sϡr�>��6���l/�{ލC���V�#�>�.i�RRO��@%ƸA���("ߥ-�J}L��8U��-�5��*q�w3O3��W�2P���̃�ִ��+�h�'n1�n{ҭ��8T�Չ�sa%Y�W���<��,�Yv������Fש�£\����WD�X!*ف�j�ǠV�:ǿ���7.�`�ƛH�0p:9[�tx���p���鏗O�4v�da���^��;���5ݎ������5Y���O�|�k_�������������t8M�C	L�l��-�^K{w7l�:ӷ��5���wG�c)�0W�]y���Ï�i]��D���LֲWU�%j��2�����͞"|KH;�oE n����t�C���g�>�Q�0ꤣȀ�[�pڗ�^>�4��?���mgd�S���x�\$�ܽs��R��3 ���K�����4D�^	�c�rԽ"8�~�lP�1�J������5�|^i�`S��Q�  9;IDAT�0&:�����|~���z�������ݑ����L&����ȅ�1W`v�7���)��7�&��v��׎����M�VG��綐�����K�`Ξ;]~�^�5>s;_��|n4$w`y��(�����%l����ľ����Óx��TƲZ��窙Z2Ԫ2Q���E�F(*-�[������ķe?�be5ߧ��p|��o� ���|~�ש�V9�ZȢܩ���,�%�K�����9�o>�T+�����w/�痮�S�,�{����'ʁ}[��"~
���i8�P��(�V����q���C�M��r��r���˽w�gh�>��wD��Tu�]�y�|��Z]_����� ��m!B��O�,w�_֠�Y~ Mg�i�7Ŏ`=y�Uj�*Ȇ��VJF]֟�������D��p�א?��!�"�Ѩ9��sZ��Pd��V�PG������UT�u��U�>�4='�.,2�v!���F�4������P�����aT� ������Y#�<�:�Q�׌���.�S�(��(N�iw9��潁B�2����j9��k!������?-���_	xK1?|�H�t�R��%C�޽s[8�e����c�� J�b��O�4����F�hP>�����X%{XV��Ӱ$M���wv�r��A-e�RӁ�)�J�K�^���qU?�Syo�>�D}M�ZQ�S�_9�Pfhf�7���7�WM%���p�:s(2Ϋ*ٵ��[�q���A!�2ǹ�@�귿������Kh��B#^oG��Lx�a�n��?���P�N �P)A��3Kt�^_E$�2-Շ�s4U�m�OS޼��/�G���f�qD�Q�����vne�me�	�|�1�q�1(�����i��5��`E9t�%5G���W#M�E��Dd�<��O}�(�rz��t3M�4�We��(�l���0��R�ݪ�QZi%�n�y"�w�̀V,M��v�kp�Ac��?"z��ܘȑtpS��!��1��O�1�4e��r� �K5�fA�B���yQ:�0xd��ԻZSR���U8J�N�5"z42��%�����H�Ը4K/�k��\�;���1��o�W��l�p�F��94��z���� �y��9�����A�ϱ�W�lq(.^�\�����!EKK�0��|f���G%e�}�m�X�A����(D���gfA'�0l��̤�%�g�h��T0�,Q5H����n� �]�3��ڊL�Ɍ�Tf��dyD�J���*w8�#�;~"�@7,&�����+o�u��/)GN�c�$��YJy�H�lr}.��w��_���L�����6��#�﾿�y��K]���2m�̿=��Se�7�](#=���������}�����o�|e�t�K�"Ѷ�M��{���i�����4V-sc\V�o��q(��-e=Zzj+�	��n�U�<TKtlz:O����c>�gk"r�K�noz��.��!hl1W!R�Ġ�J�ᘰJ9h@´�6h�>u��x>'�d!�3�N8�j2��Ʈ���J���(�wE��Q���RUG쬠a����An����*�^F�bcM��r8S�:д���^޲e�.�P�+_�V��+��;�/|����F�o~��d���K,�Za���LZ�������N�,��jo;zV8pq��]����2%G������c�Eb�!��4|{�KhJ���%�zb���2M5�QuJjQ1��ŏ�3j�V�)���q>v�n��n����!�4 q�/��`�i�����݊�%�>?Sw�o/��O�Q�8��}wc�XDw�����ʁ���W��F��Y6	*�Y"�^s��N0J|fc��
�!�N|-��S��k}��[QG&{�7ZW�(V������ ���������J��(���F��>n�V"x�U��t�v�|��("<�oȟw?�u�D]ʐ���;.�ѿ`�7;ʇ���<���[������� H.!*����ݝK7ҰH�tw,ݵt/ݰtH7�����W<�9����5��y�����̚���2��EQ���L5>���ctu^��O5�m������P'�e�e*���S�����<�9.N�.ԱQ�:tT!J����?�>|�`�r�T��&���쇴*���z�Ԗ%\��%ZeS˱7����o��^௏���;so�A�#��5�G�a�������0�**]��i���8P���%s|��9����w\:Y�+�;^�mZ�8:���kP��_����h�ޭ�y^i��K7[�/�����Y�#�Ĳ�������D�k����eѷ��p�~�L�8���iZ���hL� ѱ�����x�6���#]�4\#���p��dZ���}Z#%�Y$�)�+�r�C�,�������p�75n1Y��/0�b�p>�l?]1ׇ�S���#�lNAH�1���r��9�ԓ���P�z�zPn͟�`>���x0�;���h�����TI�~�c��c�?\�2��Z�j�.|���v?~B�N��ꃼc�g�X�`����D��&k��k�K�jW��E�d� �P�?��H�0��K�l�χ?��>���N4a��O�� �wO��]��w��jA�׷ב����PUPw�+d�KArO�cİ w��v���m���X$���3)pW&���1��u��bmC�z��6jy��{����_�� g�q���!��nh�����,|כr��|�]�yOn�ള����&i�g�(���vm��o9S��U�I��K������xN*����e����C��������S�))���_lRa'>, ���N�Ϋ�w��\�o:-�WX7\��s#��PZ>�۸N��d0�_vj2�~���=�r|��s���6��.����6��$��&ն� J<��~'�@q)줚OO��=h�.�z"�Rm㜮���R��AȟU�0�5�����+�{�r���7Rk|���h���s2�ohG�4J�\���2 ��"�)3�G��:��׬b��]A�Ň��ۭ�t/��N~X����E���#%���}�2�3_�Z�O����.�2�����M�5�
��n�5�(k��jbd ���LIf��ޞ*��XfȖw����2(�2��Jm�N����S,D%v��-�q@���j�4U�%�$�?��g�
8�s�Qo���j.�\�Z�4�^�O$�>�=뇼7�
�����}U��&�T�x
f]:Z�����8n�s���)0� �'iZ5-4ﭵ�倰,�SJ���tx�:��C4짖�O�K�+i<Ho�)�Uw?k@ן���v�ʟ�i�-�Tyފ�T*�[P�����&�t�!Eۤ ��|�o`�k"o����tJFS:m��<��4��
�����ǿ�#柕S��>����*��-����=WK�,ŞV���a�Ȗ%��s5��"�U�qQҾ-��r*e&tU���s�ӝ<j�Q�ks�7V�J�x������@��y>����R�+V�%R1$�vw_�I����1��`�_�_�|<蹩&YZ+A��d��h@�鄓����ݓwc�3�TQ{�XrRdK^8�e����?�Q�c�,����_���"�'�Iƿ��ԜΝ��G����ZfWP�Ô+�;)T@�̒�m6�$R_��d����o�;b�袜���f�v5�H2����덴��a��O0��d��O���.�P��
�|���j~a��n��v/l�~{fV	�%�!���5��;84ls�.l��5�b?�ܞ2�	�	-�VK�GٲNP��Z��熑 ���L�v�1;h�)h��K�2�T��(�7�9�ДS��:S�)�dUt�܄�m��wR@fd�+�Hs�~#�ܴ�)%�}P5|��JR��.8b;`&�j��ms����^��"�7md�A�^#��/�^�LNQ��2��A�K����`����in���x[�yCp�K����w,�s���2zgr�2QR<JZg��	��թ���:������8��r��M?�4�P�����u(L�*���!")��7Y�)b�����7�zk2@gyO����]<��&�C�<|d�|<��QuGJҬ��Zٗ��W��(G?�{��KY�F<-��8*��O�y����S�k>�u@T6c� �y�y��{OA�*�gN>��A{\i#!k%�|���X&I�61���۟ƋPZ�V�G�G�ʜ�������~��N5d�o!-�$?|]&�^�fI�ܩR�v�J�hV�(O�P����"������~�Y/�Бcߪgv0�ex�M�Bξ�@Π�[:󏺦28�;e��|��A��N�i �Ge��z�������Z>��T`�PJ�{5�x������	G�!�_�/���}@7����~�ֻ�}C�b !�	�T�raԋ��w6!��������� u��j?��[�;n��`j�;�W���+����(��Xj���o,�æ��Z����8,S���;�'��;�i�U1���g�Չ��K6���X.f_*���c!)�{��T�~Z]�Sю��S���6�S�R��ZT.���ً�PVT����� �.�T����<K�&~���q���.����V��}LR��r�DPMٞ�O9I���7�2��0��[RiE���X�x�&�й�
 ���w��?ō�M�Ҥ���Q T>Ώ�)�݄ȸ�V2|-�(�;T������+�-ڶ����?��چ������R����Ol
��/��.!���=�7�:m맵`����=Z�qkA�9�Ip䩦����{�Vm�!\j�'�:��-��S���9��	�|�v�}]���)�;�]uR��Cȵ�-�|�4���o巐������{���۹��
�ax�����p�>˜�D�G�ڽ~Y	z�u>Y����M�u�,�}Ca���wB�������Ao�־S��[dz?�跬�=��~X���jZ*#Y_�#:d	�d��w�ۀ+6�\���W��Q�O'�w{���{��am0҃){ E��No{m8�6�RͅD�޺}���D^ҫl]kφ�5�����_@�k�[�6�2��$�pxӛG��?)|��^r���_�	.x}�D`�>n)e!h��#����4l��^����|��?{�4�������s��`\��|l/��п洡�p����>�2=�Mq�``�<� (�i��E5�L����;��c�ǽ�pZZ�%�f�r�7�dҮgs�a��f=,H��{�;yg�>��Vũ�Zv^U��`�
I48Q��GڋB�)�}xU'�^7�:�Ny}y�N��s��x��M��ɋ�79JK#������lW(��jόd�}��'�
8	�����eK9+�c���Y����ֿ�q`vE�|*����M}wq��{��H��|� y�HD�X��>��^^A+kF�1j {�.[��l|�ﾊԻ��und�L�_�`%T�#��v�f�Rtl�è��9������	I=݌F�v��ʩ.\�&2�����d"m���OI#!ۃQۊ�����CN�Z���b����`'��!��ǺM|��-��%���bN�X�>�"����ciK7z�~[���_}w՘�ߔ_˔�5��{IXRV�VWV�����S���T��� 1�*)���;�N~H�-�5�wK+J�n�A�>��㳴�&�5Aë�<���^��z�ج�7k9ըM���β]��k����4,�c]��l��!f�ź�.&�%_�O�zz\敿���������`�N�gH�n�a̍v�-ܣ}^ϯ]ey�}�˴r�y�g�8Y����B4��傁p���=`���Z\����-_���o�j}G�a�����x���˯9R���S��u�X�����b^�2��C�����y���(���!+�kF���$1�ڻ���\�	Ӫ� z�����]�Ѡճ�9ۛ4<�g�5�n��?�y���L��|y&o�=�'_�T����HD�Z��ψ!����ᮾ#*H�6rZW5 �FG�	Z���Qa�w�Ӟx��.P������*ZQ�`�Z
5���y���D���aJ?����OG�'7o{�)��c渎ӂ�m�y�^YdU���R���M�S{�P�Z��-`"��z�d����g v�~��T�55����T�m�~��9:�N����xᵠE�0�wï��fb,�����%-lP�)�Rh�F�eU��a����m��\�3��vꔋ��5� �L3�;�FS�V9X�w�+Y
	IG�)3��q־����%��&�6�Xe�` �b�MK�E�?ѥ�I�?�"kg]~_���:>�C^$��vF�kx# �G�£�PI0�;.��L�?�-��ЃCF�|(X
���6C�<���]焱7��}ˬ�����-o/�1�2扰�t�����Q���Ty�<��AO��GI`��8$S��	|���!
ގ{���r]d򸤹��g�O$a	�ky��7��_��ҖFL�_���w�k1U����%���)��\�ҁT�V{Y�l�6��%x�+FJ+�eW��A�343���S�X+"�m��X��3>�	�Z�x�ͽ0/ �M���?�CF�m?S߆�L�%��c�[%�ߏ�l�����o{b�zJ��Џ�`P��9�d�po���O�"r�W7�t#l�.��������Zdi�$z�8��Y�7G[hFﰈH�s�R���	;eꜫW\����T&"�Nt�Ɩ�My��;�����	H�/q:�	��ER��^�Qרg��eU�`�|��
7j$�<���6#�Tm"��9�}�J�.��=ܓ���"��/pG�����h��耲�>j|Y���d���4N����i�a���+E��C�d�,�����	�<	Ei�+K�ym�&!Ο�)���zn�ۻ�Tf���5���L���K�}��9��H�s� \�HjM����3��6�I�]9{hW��s^��M����O�7��D�tv-���Ci�P٪b��u�gg�aH���s���(~�}�H��X*�$�cg��Y�8���QT��f��% � �TCbr��ϠVH,��ޙe��/�Gۄ����H��t"KK�R�C�����1�uϑ�Wx��i�;oؙ2%]���(jA!Q���g]|��b�)���F@!ۘ��7o>z�����xH��D)��[�����K���Ve��e��>���]��i�ƈ�~5���-��}z,]�s�+�hBw�S4h�E����IN?�Ѱ{�m����d{��듵[:xm��c��G0����7yYo�mw��� g�� �K�+'Ƭ���9�Q5,�!ȧ��Sb���rx�����.��%aM�E=�*��te�syU��"єv(�Ư�WQ���/5�u�p��T���۲��"���9��{V2�v���A��3EE#$U�+�9BOW��&fGIJO�c��
�~n�6�7]Z�&����2Wfv*$�HU����dk��U;�Ǜ�U�  �Kw<�wDe۔e�m�Hyo�0�{!B��3V&RNJ���%��l9����V��7���t�c�g����p�蒏�Aa�6��ȒRA:F;=\�1�I9:~���qK
�v���9(�25#9���HC|��G�%3�ǿ=��B��f�os[�5��J#����O9Ua�d�����5��+G����6��ظH���[�Y3��Y�8�v���k7���^\�J{����,�(>�k�C�F�nOF��k�9-'Ѓ�3�?g�,���3���3-��%'MݟD����Ӗ�7D�kj��s���Ð�f�3I�����H�H��[;�Z�˨��W�G��>NF��0-�rHq�{�L[�$��0�=��&i��)����d����E�s�x��Ӎ	�q��� �N�C����AL������ӥ��q�]��v̏o�b�@�y=�Y��?	�V�����q�J�\M��\%����_������b���4�J}�,��֍�����O7�i����(�q�Q�Yy�*�ي�9��kN����<KK��<w����P����(�"��y%r��B^'zXB��}����\}���߸�F�>`m��Nt"s�v5\��)Qv�p��6lk�PL�e�+�k)��/��:�&߽o�n��|h����m�J�rX�d�k�T9BN��$s��LU�ҷ�uAC�b	��M �b���,�y:����~,N�;�FM�����K��u�45��uތv��f�6��k�,� ��Sɵj�5O�$!�K��7���/[(Y��'��Bk��R����N'#�&�Y��	g�Axy��)����.� v*��&W���COj9�e>)�t��#|-xl*3A�R�����9:�䴹,C������l�b��6@��p�����t��l��W��k.��= ��
P䞬i��L�m+�u2������F��<�I*~�^M���R&��"�x�C�i��k}�/ST��/�mQ&�Z�K@2�elk�Qo��)���K-�i̊�P��&�������]92!�V�kЋ=�\H8��1P\"���K���������؟5�t^�;�t#e����%�q�!�&�JNhj�i����H;Y�`��
���X]��N�t�!�Ϸt3���_�Y�7"�v�[?`{
<:&1��W���_�m�Ն�m��$��<�a5K�!�e�0�}�<v�[>�%H��(-�RN�/C��������>�GEQ[��FT��S@s�Dc"�e+����%}�F��>���5�y����Mr$˫�`1..���3���.L����;�r��'dp'�X3�mK�yD_A�}-�':��Y�\�^�'��t�bb���-�x��S
���*YO!�K�
b$e�Ou?Ao��ϔӚ�n��]��JNE�'��Y���F�:���F�b̓˓�?ӳ�7�ڂ��=�fFuݑ��"{3�j륻G��̀1�?����������?\��y��|�v2�vp5�v��W�LI�����n!7� �i"�w�2�A�?ޖ'�%�/�罤%�n3��_��7��0�.<�� �t9=]��ڍ};5ZIӧ���b�d����`��X�\Q����>���q�6�<}蓚��HC�6�;�2M�*s�H%���^����}�nQ��z�F2����-Rĸ
$2C�6�5LS�C�D�2L��?CL׷���	��	)N D	�T����Z4�{u���E`#zmu��y���kP���J-oU,s{u9�s�g>I����0eu�H��;{�ڳ'K^��ߌ	���������tݰ
��X�1|��f�������#��f�6��0�Y�s���~�`����ha����E� ~��&X�EC����%0�	u�96D���j����`��k�?�٘tx2oYr8n|�q�Y�S���O<��!^���Y����ߢ�bzX=�U����{V�W�NRzp���~V�*�	�j�yj����!��Q�aE�)�B�І򖪌;( �&(���Y� �4��w��P�jog3���nOq�qI8�����ih�E�^�b.b'�ˇ,˱��fWf4�QB�|�a�0Q�Q��|���etb���*GR�ѹo�\-;-�h�0^ۚZ�>��]�-m�c�ɜ�R0I�����i�a��Hҏ,􄡬�^	_;��S�Fl=3�cg�B$��=!�����M5sg��>v.�����e�~��P<�w�X�����Ƃ�a������ꮄ��琉TQ��Nm��]����A��=�郲en�z��F�~����7�pˠZb���fʽ�H�rͨF�mE|���2MfA1�g�E�,¹�܅8�a��C\0�����w��@Z��f(�ԡC��WX�5��π����݆i� C��n��ϥA�����Z
��6�v�;#����N�%�@��g����9���.b[���5��*�������A�#�r6,���nӻ(*7eW�J�~��0���}P�9�U����M�f������}�����x��n'�<d%[��,묾F,<XZ�_;rq�����F+�v����&8t�V���__�M��^_u^ls�T<Ǡ�9�@Ӈ۝���n0h��x�D =�C�pR''N��m�<�,A�bR�k=��v����Ix6 �t�A�Ӕ�$�x�-�c���^a�t�lvEX����!3db���a^k8̒�l3J�3�l��9t؎ܯY��iŜ�Ay�zXW�<7WR��od������vB 9IX����Z�5Y?C+��p���#u���}瓊2(DR�X���r���oH)H�
�'g�d�����<h�D"���".��dw��<��vۖ�e��G��jYN-l�I�}����O�D��\�ތ�S�n�y8�[#�y����4-͝:u}�G�L�cg�yk��UM��|�٤�q�@6���/H��0Ē�?3�6B�t-Ag5��E1_t�<x�A?�v��Ot%>[ӀK��9�U�¤m�u�Y���{��uI�hGH�[�UH4D�Ai:M���̕��A� a���.�?�?�h�FgKu�M��վ g$�J��gѧ�e���|?���=��|���<PB�r��R8�֥sI���ZKV����:t�R]��D���_�]Y����0ڍ�Cg�F�ը��9�V9e�r�^�{��3e���H��(Jw<\h��Q��M2F?<�0?SV���>7/�Pg-zB�$�:/=���i�{Z�ХO.�{��R5��ۭ�!�aR�U%��3���C|�z���A��^}����OSq1Iy�ki�����_�i��<�Gu~ZP �'��f]�I�N��͸̏!w�M����b�ߗ�"�)��-��A~R�Y�����6���dZ������o��Uc!���@��Dx��s��у�"k`�w�Դv��F{������Sj�r,���Z� -�������fO{�e�7�F��ܢ]&��;���@�7w�%cԆ����3�wv�Ļ.:s�����>η�x+�m�p��a��}6r�Xy�V���~�S�#��2��`��e�I� I$ڣR��`V	`t��xŔ+��Eg`���nf�6��Aa�W(C����
��^h[�2����f֐$k����[r3,���>*�U	a���6��G}+�J��
�n;8�Tp#�U��E��PIT�0W�֨�b͛�C��]}�?<*{�R�U�v�˺�]�^q=kf��#�c�wB+�|�o1�߉���0��ܫ��Y%hOMH�cO���� �D���W�ʝA���+8Kp�k�u�nG�.��#�{Y��s��y��A9��������N8�O�'�XP��˼��V� ���J�)���Nj�2VJ�Q��Y&��f���� �)��+�' p�LK�-��h�T�3�>��"�3��R�aЏ��b=6v��k�0�W*����}�J	����]䯯Y�J��3l��i(3�����]�4�}��pߤ�!�I�GG��JJ�
��N��2�o�hwf����Ѷ&���)�޾���"�]�#ɹ��+�3��+��'+e^�.���]�\H[�g�ʝ�Ck(I+��K���������>�F�b8P�<�=�ݜ'�ĕ�M��p�o�-�M�Ӄ�~7��F�ܩ+R]�ﰾ۟��r�=��s�Y��W�=�r�'�Ǩ�s(���H@�Oҳ���(W�ͼ� �޵��M=�Wn�F���Q;��yۥ.�"6Ih����J?Ȁ
����fq���SŌ�d<+ۡ8*KϠ~H�����@���4�^a�;���	��ZcҺ̠��dM�˙g�`K�co/���Pc�ץEԤ�3���:YVOa��� ����JJj�}��/ɭ2�	Jx�fv��M��Quu��]�eǮ#$��d���2)���%�X�F~���%�[�Ѡ����k��͐�9�-�&T�dlʌ�]*I�$`.g_��1MiP��[�ݧ�P�*JD$7��o��8� ޏ���;�ߴ+9�����^��o����l��# ��R��x+N�����>�̾�q7G��y�H�����ޕ�g��}WD���GIPT&(uM�Dk�����Zw�p�byz����"/R��l��}'	17�M�=#�oo9爑�<%��mIl��y��Vm��\�z���XU��&�@�����ȁu��W����*4)r�[R1���t�i#�W�K2f���E�u���+�"�g�8�!z& ���ƮZ�?ʠ�9�,m՞��˓���u��L��$N���J�V79=��gm��l�%4�.�^K:����g�����B���:�\�����$l雼�^8��{/��15��Y�d�%�B���c?tI��u��*mrx���\��Q�<Et~��FSLa�b&d`�\4Q���6V-��� �I���s�Oz[�u�E{�㼡�6|�@�nH�z'_�OU׷�4�6�5�"؞X^8ǐ0����f����&���Q W׌{�۴9܇d�a�v�v��>����_��1oY\_s!zYȟn�6����BϷƆq�7Dwe�G�-�PQ��nKk�|����$�ݾ����0:r�y�P�a�7�3��I<�"��bح�g�������^�h���`�CoV�t���X�,�:`��烼�t��2�dX���5:��(�r)�����x�6M˔i�G���ҏF}�,�R�^�����|�j�t��<����t�|:���-Xb��j���q����y�C9�fv�Ys�ď]xbS�l�X7>�m ���A:�"���T"�f�� �z�8
�˶/&���=|�{�bY���<<�s�p�T���V_��(��s���s&��5��Q�\����v>^��wMq���>O���-:�^�o��,�z�ͺ���j����a���突��cJ�i���5� �<3�sku�W���rU�Q5�}�=�:,t��[L�p�tXv9j}��:�:�������?�����?��	Yj�/���1=6��o�3IE�J1���PK   ?To���!       jsons/user_defined.json��;O�0��
�\[vb�IV�0� ��*�*K�9	UU�s�]:�l�s�9��߷�h�l�4��`Z�/�:(���K7�Iڡ��p�<5�i��KP覷���@�`w�<ۭ��i�������s�d��Bb�U�*��S�T�Z�i�?�K�������Z�����k�k}x.���°]���4�����!V^RY��:{���"2�<YL,V���	��'�<�S��M��g��1��丸�9��YUJ@�Ì��h���W�p�*���9�s0Rf�ɛ�)����1�.9��oPK
   ?T$�2@'  �~                  cirkitFile.jsonPK
   /�>T�a��V _ /             m'  images/b9b5db0f-1139-4dc1-aec6-3976f40bff5b.pngPK
   U�>T|p - �9 /             �~ images/cdb0e0ab-4d76-4fa2-8457-7cb33d05bd01.pngPK
   ?To���!                 � jsons/user_defined.jsonPK      <  <�   